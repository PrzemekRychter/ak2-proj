* NGSPICE file created from adder.ext - technology: scmos

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt adder gnd vdd S[5] S[4] S[3] S[2] S[1] S[0] X[5] X[4] X[3] X[2] X[1] X[0]
+ Y[5] Y[4] Y[3] Y[2] Y[1] Y[0] cout
X_66_ Y[0] gnd _64_/A vdd INVX1
XSFILL1880x2050 gnd vdd FILL
X_49_ _49_/A gnd _49_/Y vdd INVX1
X_83_ _86_/Y _82_/Y gnd _49_/A vdd NOR2X1
X_65_ Y[0] X[0] gnd _65_/Y vdd XOR2X1
X_82_ X[4] gnd _82_/Y vdd INVX1
XSFILL4840x1050 gnd vdd FILL
X_48_ _46_/Y _47_/Y gnd _31_/A vdd NAND2X1
X_81_ Y[3] gnd _78_/A vdd INVX1
X_63_ X[0] gnd _64_/B vdd INVX1
X_64_ _64_/A _64_/B gnd _64_/Y vdd NOR2X1
X_47_ _47_/A _58_/Y gnd _47_/Y vdd NAND2X1
X_80_ Y[3] X[3] gnd _80_/Y vdd XOR2X1
XFILL5880x2050 gnd vdd FILL
X_62_ _62_/A _50_/B gnd _53_/B vdd AND2X2
X_46_ _57_/Y gnd _46_/Y vdd INVX1
X_29_ _47_/A _29_/B gnd _35_/A vdd XOR2X1
X_28_ _64_/Y _70_/Y gnd _28_/Y vdd XOR2X1
X_61_ _61_/A _61_/B gnd _52_/A vdd NAND2X1
X_45_ _45_/A _44_/Y gnd _45_/Y vdd NAND2X1
X_44_ _47_/A _74_/Y gnd _44_/Y vdd NAND2X1
XSFILL4760x50 gnd vdd FILL
X_60_ _49_/A _62_/A gnd _61_/B vdd NAND2X1
X_43_ _56_/A gnd _45_/A vdd INVX1
XSFILL1640x50 gnd vdd FILL
X_42_ _42_/A _42_/B gnd _47_/A vdd NAND2X1
X_41_ _64_/Y _69_/Y gnd _42_/B vdd NAND2X1
XFILL5800x50 gnd vdd FILL
XSFILL1960x2050 gnd vdd FILL
X_40_ _68_/Y gnd _42_/A vdd INVX1
XSFILL1800x2050 gnd vdd FILL
X_79_ _78_/A _78_/B gnd _56_/B vdd NAND2X1
X_78_ _78_/A _78_/B gnd _78_/Y vdd NOR2X1
X_77_ X[3] gnd _78_/B vdd INVX1
X_76_ Y[2] gnd _73_/A vdd INVX1
XSFILL4840x50 gnd vdd FILL
X_59_ _59_/A gnd _61_/A vdd INVX1
X_58_ _56_/B _74_/Y gnd _58_/Y vdd AND2X2
XSFILL1640x1050 gnd vdd FILL
X_75_ Y[2] X[2] gnd _29_/B vdd XOR2X1
X_91_ Y[5] gnd _91_/Y vdd INVX1
X_57_ _55_/Y _56_/Y gnd _57_/Y vdd NAND2X1
X_74_ _73_/A _73_/B gnd _74_/Y vdd NAND2X1
X_90_ Y[5] X[5] gnd _90_/Y vdd XOR2X1
XSFILL4680x1050 gnd vdd FILL
X_39_ _39_/A gnd cout vdd BUFX2
X_56_ _56_/A _56_/B gnd _56_/Y vdd NAND2X1
X_73_ _73_/A _73_/B gnd _56_/A vdd NOR2X1
X_38_ _32_/Y gnd S[5] vdd BUFX2
XSFILL5080x2050 gnd vdd FILL
X_55_ _78_/Y gnd _55_/Y vdd INVX1
X_72_ X[2] gnd _73_/B vdd INVX1
X_37_ _31_/Y gnd S[4] vdd BUFX2
X_71_ Y[1] gnd _69_/A vdd INVX1
X_54_ _54_/A _54_/B gnd _39_/A vdd NAND2X1
XSFILL1480x50 gnd vdd FILL
XSFILL4920x2050 gnd vdd FILL
X_70_ Y[1] X[1] gnd _70_/Y vdd XOR2X1
X_53_ _31_/A _53_/B gnd _54_/B vdd NAND2X1
X_36_ _30_/Y gnd S[3] vdd BUFX2
X_52_ _52_/A gnd _54_/A vdd INVX1
X_35_ _35_/A gnd S[2] vdd BUFX2
X_34_ _28_/Y gnd S[1] vdd BUFX2
X_51_ _49_/Y _51_/B gnd _51_/Y vdd NAND2X1
XSFILL1720x1050 gnd vdd FILL
X_33_ _65_/Y gnd S[0] vdd BUFX2
X_50_ _31_/A _50_/B gnd _51_/B vdd NAND2X1
X_32_ _51_/Y _90_/Y gnd _32_/Y vdd XOR2X1
XFILL5880x50 gnd vdd FILL
X_31_ _31_/A _85_/Y gnd _31_/Y vdd XOR2X1
XSFILL4760x1050 gnd vdd FILL
X_30_ _45_/Y _80_/Y gnd _30_/Y vdd XOR2X1
X_89_ _91_/Y _87_/Y gnd _62_/A vdd NAND2X1
XSFILL5000x2050 gnd vdd FILL
X_88_ _91_/Y _87_/Y gnd _59_/A vdd NOR2X1
X_87_ X[5] gnd _87_/Y vdd INVX1
XSFILL4680x50 gnd vdd FILL
XSFILL1560x50 gnd vdd FILL
X_69_ _69_/A _69_/B gnd _69_/Y vdd NAND2X1
X_86_ Y[4] gnd _86_/Y vdd INVX1
X_68_ _69_/A _69_/B gnd _68_/Y vdd NOR2X1
X_85_ Y[4] X[4] gnd _85_/Y vdd XOR2X1
XSFILL1800x1050 gnd vdd FILL
X_67_ X[1] gnd _69_/B vdd INVX1
X_84_ _86_/Y _82_/Y gnd _50_/B vdd NAND2X1
.ends

