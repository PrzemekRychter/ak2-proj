magic
tech scmos
timestamp 1590258663
<< metal1 >>
rect 469 307 475 308
rect 464 303 465 307
rect 469 303 470 307
rect 474 303 475 307
rect 479 303 480 307
rect 469 302 475 303
rect 78 271 81 278
rect 118 271 121 281
rect 70 268 81 271
rect 102 268 121 271
rect 194 268 209 271
rect 254 262 257 271
rect 530 268 537 271
rect 86 258 94 261
rect 142 258 161 261
rect 302 261 305 268
rect 302 258 313 261
rect 394 258 401 261
rect 158 248 161 258
rect 233 248 238 252
rect 561 248 566 252
rect 426 238 433 241
rect 630 238 646 241
rect 506 218 521 221
rect 173 207 179 208
rect 168 203 169 207
rect 173 203 174 207
rect 178 203 179 207
rect 183 203 184 207
rect 173 202 179 203
rect 298 168 305 171
rect 94 161 97 168
rect 414 166 418 168
rect 86 158 97 161
rect 274 158 281 161
rect 214 148 249 151
rect 558 151 561 161
rect 558 148 577 151
rect 58 138 65 141
rect 138 138 145 141
rect 162 138 193 141
rect 318 138 337 141
rect 342 138 361 141
rect 366 138 377 141
rect 382 138 398 141
rect 442 138 449 141
rect 582 141 585 148
rect 534 138 545 141
rect 582 138 593 141
rect 62 128 65 138
rect 126 128 134 131
rect 358 128 361 138
rect 410 118 411 122
rect 469 107 475 108
rect 464 103 465 107
rect 469 103 470 107
rect 474 103 475 107
rect 479 103 480 107
rect 469 102 475 103
rect 78 68 86 71
rect 126 68 137 71
rect 398 71 401 81
rect 382 68 393 71
rect 398 68 417 71
rect 422 68 433 71
rect 462 68 518 71
rect 622 68 646 71
rect 22 58 57 61
rect 94 58 113 61
rect 110 48 113 58
rect 358 58 377 61
rect 510 58 521 61
rect 554 58 561 61
rect 246 51 249 58
rect 518 52 521 58
rect 238 48 249 51
rect 454 48 462 51
rect 534 48 545 51
rect 534 42 537 48
rect 173 7 179 8
rect 168 3 169 7
rect 173 3 174 7
rect 178 3 179 7
rect 183 3 184 7
rect 173 2 179 3
<< m2contact >>
rect 460 303 464 307
rect 465 303 469 307
rect 470 303 474 307
rect 475 303 479 307
rect 480 303 484 307
rect 278 288 282 292
rect 414 288 418 292
rect 606 288 610 292
rect 6 278 10 282
rect 78 278 82 282
rect 110 278 114 282
rect 14 268 18 272
rect 22 268 26 272
rect 302 278 306 282
rect 318 278 322 282
rect 326 278 330 282
rect 334 278 338 282
rect 422 278 426 282
rect 526 278 530 282
rect 134 268 138 272
rect 174 268 178 272
rect 190 268 194 272
rect 294 268 298 272
rect 302 268 306 272
rect 342 268 346 272
rect 390 268 394 272
rect 438 268 442 272
rect 486 268 490 272
rect 526 268 530 272
rect 582 268 586 272
rect 46 258 50 262
rect 94 258 98 262
rect 254 258 258 262
rect 262 258 266 262
rect 286 258 290 262
rect 366 258 370 262
rect 390 258 394 262
rect 462 258 466 262
rect 590 258 594 262
rect 614 258 618 262
rect 150 248 154 252
rect 238 248 242 252
rect 566 248 570 252
rect 422 238 426 242
rect 646 238 650 242
rect 126 218 130 222
rect 166 218 170 222
rect 502 218 506 222
rect 164 203 168 207
rect 169 203 173 207
rect 174 203 178 207
rect 179 203 183 207
rect 184 203 188 207
rect 262 188 266 192
rect 550 188 554 192
rect 614 188 618 192
rect 94 168 98 172
rect 294 168 298 172
rect 414 168 418 172
rect 494 168 498 172
rect 110 158 114 162
rect 158 158 162 162
rect 270 158 274 162
rect 286 158 290 162
rect 310 158 314 162
rect 350 158 354 162
rect 390 158 394 162
rect 462 158 466 162
rect 70 148 74 152
rect 134 148 138 152
rect 438 148 442 152
rect 510 148 514 152
rect 566 158 570 162
rect 582 148 586 152
rect 6 138 10 142
rect 54 138 58 142
rect 94 138 98 142
rect 134 138 138 142
rect 158 138 162 142
rect 238 138 242 142
rect 270 138 274 142
rect 294 138 298 142
rect 398 138 402 142
rect 438 138 442 142
rect 518 138 522 142
rect 638 138 642 142
rect 78 128 82 132
rect 102 128 106 132
rect 118 128 122 132
rect 134 128 138 132
rect 150 128 154 132
rect 326 128 330 132
rect 422 128 426 132
rect 454 128 458 132
rect 526 128 530 132
rect 30 118 34 122
rect 406 118 410 122
rect 430 118 434 122
rect 460 103 464 107
rect 465 103 469 107
rect 470 103 474 107
rect 475 103 479 107
rect 480 103 484 107
rect 110 88 114 92
rect 198 88 202 92
rect 286 88 290 92
rect 310 88 314 92
rect 326 88 330 92
rect 518 88 522 92
rect 598 88 602 92
rect 142 78 146 82
rect 230 78 234 82
rect 246 78 250 82
rect 318 78 322 82
rect 30 68 34 72
rect 86 68 90 72
rect 174 68 178 72
rect 222 68 226 72
rect 254 68 258 72
rect 262 68 266 72
rect 294 68 298 72
rect 438 78 442 82
rect 494 78 498 82
rect 550 78 554 82
rect 566 78 570 82
rect 518 68 522 72
rect 534 68 538 72
rect 574 68 578 72
rect 646 68 650 72
rect 102 48 106 52
rect 246 58 250 62
rect 270 58 274 62
rect 334 58 338 62
rect 550 58 554 62
rect 310 48 314 52
rect 366 48 370 52
rect 406 48 410 52
rect 446 48 450 52
rect 462 48 466 52
rect 518 48 522 52
rect 6 38 10 42
rect 534 38 538 42
rect 342 18 346 22
rect 164 3 168 7
rect 169 3 173 7
rect 174 3 178 7
rect 179 3 183 7
rect 184 3 188 7
<< metal2 >>
rect 78 338 82 342
rect 254 338 258 342
rect 270 341 274 342
rect 270 338 281 341
rect 78 282 81 338
rect 254 312 257 338
rect 278 292 281 338
rect 318 338 322 342
rect 342 338 346 342
rect 406 341 410 342
rect 406 338 417 341
rect 318 282 321 338
rect 342 312 345 338
rect 334 308 342 311
rect 326 282 329 288
rect 334 282 337 308
rect 306 278 310 281
rect 6 252 9 278
rect 14 272 17 278
rect 110 272 113 278
rect 318 272 321 278
rect 390 272 393 308
rect 414 292 417 338
rect 438 338 442 342
rect 518 341 522 342
rect 598 341 602 342
rect 518 338 529 341
rect 598 338 609 341
rect 438 282 441 338
rect 469 307 475 308
rect 464 303 465 307
rect 469 303 470 307
rect 474 303 475 307
rect 479 303 480 307
rect 469 302 475 303
rect 526 282 529 338
rect 606 292 609 338
rect 426 278 430 281
rect 438 272 441 278
rect 486 272 489 278
rect 130 268 134 271
rect 178 268 182 271
rect 290 268 294 271
rect 338 268 342 271
rect 22 252 25 268
rect 190 262 193 268
rect 254 262 257 268
rect 302 262 305 268
rect 526 262 529 268
rect 50 258 54 261
rect 290 258 294 261
rect 362 258 366 261
rect 394 258 398 261
rect 466 258 470 261
rect 94 252 97 258
rect 262 252 265 258
rect 146 248 150 251
rect 234 248 238 251
rect 562 248 566 251
rect 166 222 169 228
rect 94 162 97 168
rect 106 158 110 161
rect 6 142 9 148
rect 54 142 57 158
rect 74 148 78 151
rect 94 142 97 148
rect 98 138 102 141
rect 126 141 129 218
rect 150 161 153 218
rect 173 207 179 208
rect 168 203 169 207
rect 173 203 174 207
rect 178 203 179 207
rect 183 203 184 207
rect 173 202 179 203
rect 262 192 265 238
rect 298 168 302 171
rect 350 162 353 168
rect 414 162 417 168
rect 150 158 158 161
rect 274 158 278 161
rect 386 158 390 161
rect 134 152 137 158
rect 126 138 134 141
rect 78 132 81 138
rect 118 132 121 138
rect 142 131 145 138
rect 138 128 145 131
rect 30 72 33 118
rect 86 72 89 118
rect 102 62 105 128
rect 110 92 113 108
rect 142 82 145 128
rect 150 122 153 128
rect 158 112 161 138
rect 238 92 241 138
rect 270 122 273 138
rect 286 92 289 158
rect 294 132 297 138
rect 310 92 313 158
rect 402 138 406 141
rect 422 132 425 238
rect 490 168 494 171
rect 502 162 505 218
rect 582 192 585 268
rect 590 252 593 258
rect 614 192 617 258
rect 646 242 649 248
rect 554 188 558 191
rect 466 158 470 161
rect 438 152 441 158
rect 566 152 569 158
rect 514 148 518 151
rect 438 132 441 138
rect 446 128 454 131
rect 326 92 329 128
rect 434 118 441 121
rect 202 88 206 91
rect 310 82 313 88
rect 242 78 246 81
rect 174 72 177 78
rect 222 72 225 78
rect 230 72 233 78
rect 262 72 265 78
rect 318 72 321 78
rect 250 68 254 71
rect 298 68 302 71
rect 102 52 105 58
rect 6 42 9 48
rect 174 22 177 68
rect 173 7 179 8
rect 168 3 169 7
rect 173 3 174 7
rect 178 3 179 7
rect 183 3 184 7
rect 173 2 179 3
rect 198 -18 201 18
rect 198 -22 202 -18
rect 214 -19 218 -18
rect 222 -19 225 68
rect 406 62 409 118
rect 438 82 441 118
rect 266 58 270 61
rect 246 52 249 58
rect 334 52 337 58
rect 366 52 369 58
rect 446 52 449 128
rect 469 107 475 108
rect 464 103 465 107
rect 469 103 470 107
rect 474 103 475 107
rect 479 103 480 107
rect 469 102 475 103
rect 510 91 513 148
rect 582 142 585 148
rect 518 132 521 138
rect 510 88 518 91
rect 526 81 529 128
rect 638 92 641 138
rect 602 88 606 91
rect 518 78 529 81
rect 562 78 566 81
rect 494 72 497 78
rect 518 72 521 78
rect 550 72 553 78
rect 646 72 649 78
rect 530 68 534 71
rect 570 68 574 71
rect 534 62 537 68
rect 546 58 550 61
rect 306 48 310 51
rect 410 48 414 51
rect 458 48 462 51
rect 522 48 526 51
rect 534 42 537 48
rect 214 -22 225 -19
rect 342 -19 345 18
rect 574 -18 577 68
rect 646 52 649 68
rect 350 -19 354 -18
rect 342 -22 354 -19
rect 574 -22 578 -18
<< m3contact >>
rect 254 308 258 312
rect 342 308 346 312
rect 390 308 394 312
rect 326 288 330 292
rect 14 278 18 282
rect 310 278 314 282
rect 460 303 464 307
rect 465 303 469 307
rect 470 303 474 307
rect 475 303 479 307
rect 480 303 484 307
rect 430 278 434 282
rect 438 278 442 282
rect 486 278 490 282
rect 526 278 530 282
rect 110 268 114 272
rect 126 268 130 272
rect 182 268 186 272
rect 254 268 258 272
rect 286 268 290 272
rect 318 268 322 272
rect 334 268 338 272
rect 54 258 58 262
rect 190 258 194 262
rect 294 258 298 262
rect 302 258 306 262
rect 358 258 362 262
rect 398 258 402 262
rect 470 258 474 262
rect 526 258 530 262
rect 6 248 10 252
rect 22 248 26 252
rect 94 248 98 252
rect 142 248 146 252
rect 230 248 234 252
rect 262 248 266 252
rect 558 248 562 252
rect 262 238 266 242
rect 166 228 170 232
rect 150 218 154 222
rect 54 158 58 162
rect 94 158 98 162
rect 102 158 106 162
rect 6 148 10 152
rect 78 148 82 152
rect 94 148 98 152
rect 78 138 82 142
rect 102 138 106 142
rect 118 138 122 142
rect 134 158 138 162
rect 164 203 168 207
rect 169 203 173 207
rect 174 203 178 207
rect 179 203 183 207
rect 184 203 188 207
rect 302 168 306 172
rect 350 168 354 172
rect 278 158 282 162
rect 382 158 386 162
rect 414 158 418 162
rect 142 138 146 142
rect 86 118 90 122
rect 110 108 114 112
rect 150 118 154 122
rect 158 108 162 112
rect 270 118 274 122
rect 294 128 298 132
rect 406 138 410 142
rect 486 168 490 172
rect 590 248 594 252
rect 646 248 650 252
rect 558 188 562 192
rect 582 188 586 192
rect 438 158 442 162
rect 470 158 474 162
rect 502 158 506 162
rect 518 148 522 152
rect 566 148 570 152
rect 422 128 426 132
rect 438 128 442 132
rect 454 128 458 132
rect 206 88 210 92
rect 238 88 242 92
rect 174 78 178 82
rect 222 78 226 82
rect 238 78 242 82
rect 262 78 266 82
rect 310 78 314 82
rect 230 68 234 72
rect 246 68 250 72
rect 302 68 306 72
rect 318 68 322 72
rect 102 58 106 62
rect 6 48 10 52
rect 174 18 178 22
rect 198 18 202 22
rect 164 3 168 7
rect 169 3 173 7
rect 174 3 178 7
rect 179 3 183 7
rect 184 3 188 7
rect 262 58 266 62
rect 366 58 370 62
rect 406 58 410 62
rect 460 103 464 107
rect 465 103 469 107
rect 470 103 474 107
rect 475 103 479 107
rect 480 103 484 107
rect 582 138 586 142
rect 518 128 522 132
rect 606 88 610 92
rect 638 88 642 92
rect 558 78 562 82
rect 646 78 650 82
rect 494 68 498 72
rect 526 68 530 72
rect 550 68 554 72
rect 566 68 570 72
rect 534 58 538 62
rect 542 58 546 62
rect 246 48 250 52
rect 302 48 306 52
rect 334 48 338 52
rect 414 48 418 52
rect 454 48 458 52
rect 526 48 530 52
rect 534 48 538 52
rect 646 48 650 52
<< metal3 >>
rect 258 308 262 311
rect 346 308 390 311
rect 469 307 475 308
rect 469 302 475 303
rect 302 278 310 281
rect 326 281 329 288
rect 314 278 329 281
rect 434 278 438 281
rect 490 278 526 281
rect 14 271 17 278
rect 14 268 110 271
rect 114 268 126 271
rect 186 268 254 271
rect 258 268 286 271
rect 322 268 334 271
rect 58 258 190 261
rect 298 258 302 261
rect 362 258 398 261
rect 474 258 526 261
rect -26 251 -22 252
rect -26 248 6 251
rect 10 248 22 251
rect 98 248 142 251
rect 234 248 262 251
rect 562 248 590 251
rect 670 251 674 252
rect 650 248 674 251
rect 258 238 262 241
rect 166 221 169 228
rect 154 218 169 221
rect 173 207 179 208
rect 173 202 179 203
rect 562 188 582 191
rect 306 168 350 171
rect 414 168 486 171
rect 414 162 417 168
rect -26 161 -22 162
rect -26 158 54 161
rect 98 158 102 161
rect 106 158 134 161
rect 282 158 382 161
rect 442 158 470 161
rect 474 158 502 161
rect 82 148 94 151
rect 522 148 566 151
rect -26 141 -22 142
rect 6 141 9 148
rect -26 138 78 141
rect 106 138 118 141
rect 146 138 297 141
rect 410 138 582 141
rect 294 132 297 138
rect 426 128 438 131
rect 458 128 518 131
rect 90 118 150 121
rect 154 118 270 121
rect 114 108 158 111
rect 469 107 475 108
rect 469 102 475 103
rect 210 88 238 91
rect 610 88 638 91
rect 226 78 238 81
rect 266 78 310 81
rect 562 78 646 81
rect 174 71 177 78
rect 174 68 230 71
rect 250 68 302 71
rect 306 68 318 71
rect 498 68 526 71
rect 554 68 566 71
rect 106 58 262 61
rect 370 58 406 61
rect 538 58 542 61
rect -26 51 -22 52
rect -26 48 6 51
rect 250 48 302 51
rect 306 48 334 51
rect 418 48 454 51
rect 530 48 534 51
rect 670 51 674 52
rect 650 48 674 51
rect 178 18 198 21
rect 173 7 179 8
rect 173 2 179 3
<< m4contact >>
rect 262 308 266 312
rect 461 303 464 307
rect 464 303 465 307
rect 467 303 469 307
rect 469 303 470 307
rect 470 303 471 307
rect 473 303 474 307
rect 474 303 475 307
rect 475 303 477 307
rect 479 303 480 307
rect 480 303 483 307
rect 254 238 258 242
rect 165 203 168 207
rect 168 203 169 207
rect 171 203 173 207
rect 173 203 174 207
rect 174 203 175 207
rect 177 203 178 207
rect 178 203 179 207
rect 179 203 181 207
rect 183 203 184 207
rect 184 203 187 207
rect 461 103 464 107
rect 464 103 465 107
rect 467 103 469 107
rect 469 103 470 107
rect 470 103 471 107
rect 473 103 474 107
rect 474 103 475 107
rect 475 103 477 107
rect 479 103 480 107
rect 480 103 483 107
rect 165 3 168 7
rect 168 3 169 7
rect 171 3 173 7
rect 173 3 174 7
rect 174 3 175 7
rect 177 3 178 7
rect 178 3 179 7
rect 179 3 181 7
rect 183 3 184 7
rect 184 3 187 7
<< metal4 >>
rect 254 308 262 311
rect 254 242 257 308
rect 469 307 475 308
rect 469 302 475 303
rect 173 207 179 208
rect 173 202 179 203
rect 469 107 475 108
rect 469 102 475 103
rect 173 7 179 8
rect 173 2 179 3
<< m5contact >>
rect 460 303 461 307
rect 461 303 464 307
rect 465 303 467 307
rect 467 303 469 307
rect 470 303 471 307
rect 471 303 473 307
rect 473 303 474 307
rect 475 303 477 307
rect 477 303 479 307
rect 480 303 483 307
rect 483 303 484 307
rect 164 203 165 207
rect 165 203 168 207
rect 169 203 171 207
rect 171 203 173 207
rect 174 203 175 207
rect 175 203 177 207
rect 177 203 178 207
rect 179 203 181 207
rect 181 203 183 207
rect 184 203 187 207
rect 187 203 188 207
rect 460 103 461 107
rect 461 103 464 107
rect 465 103 467 107
rect 467 103 469 107
rect 470 103 471 107
rect 471 103 473 107
rect 473 103 474 107
rect 475 103 477 107
rect 477 103 479 107
rect 480 103 483 107
rect 483 103 484 107
rect 164 3 165 7
rect 165 3 168 7
rect 169 3 171 7
rect 171 3 173 7
rect 174 3 175 7
rect 175 3 177 7
rect 177 3 178 7
rect 179 3 181 7
rect 181 3 183 7
rect 184 3 187 7
rect 187 3 188 7
<< metal5 >>
rect 469 307 475 308
rect 464 303 465 307
rect 479 303 480 307
rect 471 302 473 303
rect 173 207 179 208
rect 168 203 169 207
rect 183 203 184 207
rect 175 202 177 203
rect 469 107 475 108
rect 464 103 465 107
rect 479 103 480 107
rect 471 102 473 103
rect 173 7 179 8
rect 168 3 169 7
rect 183 3 184 7
rect 175 2 177 3
<< m6contact >>
rect 466 303 469 307
rect 469 303 470 307
rect 470 303 471 307
rect 473 303 474 307
rect 474 303 475 307
rect 475 303 478 307
rect 466 302 471 303
rect 473 302 478 303
rect 170 203 173 207
rect 173 203 174 207
rect 174 203 175 207
rect 177 203 178 207
rect 178 203 179 207
rect 179 203 182 207
rect 170 202 175 203
rect 177 202 182 203
rect 466 103 469 107
rect 469 103 470 107
rect 470 103 471 107
rect 473 103 474 107
rect 474 103 475 107
rect 475 103 478 107
rect 466 102 471 103
rect 473 102 478 103
rect 170 3 173 7
rect 173 3 174 7
rect 174 3 175 7
rect 177 3 178 7
rect 178 3 179 7
rect 179 3 182 7
rect 170 2 175 3
rect 177 2 182 3
<< metal6 >>
rect 164 207 188 307
rect 164 202 170 207
rect 175 202 177 207
rect 182 202 188 207
rect 164 7 188 202
rect 164 2 170 7
rect 175 2 177 7
rect 182 2 188 7
rect 164 -6 188 2
rect 460 302 466 307
rect 471 302 473 307
rect 478 302 484 307
rect 460 107 484 302
rect 460 102 466 107
rect 471 102 473 107
rect 478 102 484 107
rect 460 -6 484 102
use BUFX2  _35_
timestamp 1590258663
transform -1 0 28 0 -1 105
box -2 -3 26 103
use XOR2X1  _29_
timestamp 1590258663
transform -1 0 84 0 -1 105
box -2 -3 58 103
use XOR2X1  _75_
timestamp 1590258663
transform -1 0 60 0 1 105
box -2 -3 58 103
use INVX1  _76_
timestamp 1590258663
transform 1 0 60 0 1 105
box -2 -3 18 103
use NAND2X1  _44_
timestamp 1590258663
transform 1 0 84 0 -1 105
box -2 -3 26 103
use NAND2X1  _45_
timestamp 1590258663
transform -1 0 132 0 -1 105
box -2 -3 26 103
use INVX1  _72_
timestamp 1590258663
transform 1 0 76 0 1 105
box -2 -3 18 103
use NAND2X1  _74_
timestamp 1590258663
transform 1 0 92 0 1 105
box -2 -3 26 103
use NOR2X1  _73_
timestamp 1590258663
transform 1 0 116 0 1 105
box -2 -3 26 103
use INVX1  _43_
timestamp 1590258663
transform -1 0 148 0 -1 105
box -2 -3 18 103
use XOR2X1  _80_
timestamp 1590258663
transform -1 0 228 0 -1 105
box -2 -3 58 103
use NAND2X1  _42_
timestamp 1590258663
transform 1 0 140 0 1 105
box -2 -3 26 103
use FILL  SFILL1480x50
timestamp 1590258663
transform -1 0 156 0 -1 105
box -2 -3 10 103
use FILL  SFILL1560x50
timestamp 1590258663
transform -1 0 164 0 -1 105
box -2 -3 10 103
use FILL  SFILL1640x50
timestamp 1590258663
transform -1 0 172 0 -1 105
box -2 -3 10 103
use FILL  SFILL1640x1050
timestamp 1590258663
transform 1 0 164 0 1 105
box -2 -3 10 103
use FILL  SFILL1720x1050
timestamp 1590258663
transform 1 0 172 0 1 105
box -2 -3 10 103
use FILL  SFILL1800x1050
timestamp 1590258663
transform 1 0 180 0 1 105
box -2 -3 10 103
use INVX1  _77_
timestamp 1590258663
transform 1 0 228 0 -1 105
box -2 -3 18 103
use INVX1  _81_
timestamp 1590258663
transform 1 0 244 0 -1 105
box -2 -3 18 103
use XOR2X1  _30_
timestamp 1590258663
transform 1 0 188 0 1 105
box -2 -3 58 103
use BUFX2  _36_
timestamp 1590258663
transform 1 0 244 0 1 105
box -2 -3 26 103
use AND2X2  _58_
timestamp 1590258663
transform 1 0 260 0 -1 105
box -2 -3 34 103
use NAND2X1  _79_
timestamp 1590258663
transform 1 0 292 0 -1 105
box -2 -3 26 103
use NAND2X1  _47_
timestamp 1590258663
transform 1 0 268 0 1 105
box -2 -3 26 103
use NAND2X1  _56_
timestamp 1590258663
transform 1 0 292 0 1 105
box -2 -3 26 103
use NOR2X1  _78_
timestamp 1590258663
transform 1 0 316 0 -1 105
box -2 -3 26 103
use BUFX2  _39_
timestamp 1590258663
transform -1 0 364 0 -1 105
box -2 -3 26 103
use NAND2X1  _54_
timestamp 1590258663
transform -1 0 388 0 -1 105
box -2 -3 26 103
use INVX1  _55_
timestamp 1590258663
transform -1 0 332 0 1 105
box -2 -3 18 103
use NAND2X1  _57_
timestamp 1590258663
transform 1 0 332 0 1 105
box -2 -3 26 103
use INVX1  _46_
timestamp 1590258663
transform 1 0 356 0 1 105
box -2 -3 18 103
use INVX1  _52_
timestamp 1590258663
transform -1 0 404 0 -1 105
box -2 -3 18 103
use NAND2X1  _61_
timestamp 1590258663
transform -1 0 428 0 -1 105
box -2 -3 26 103
use INVX1  _59_
timestamp 1590258663
transform -1 0 444 0 -1 105
box -2 -3 18 103
use NAND2X1  _48_
timestamp 1590258663
transform 1 0 372 0 1 105
box -2 -3 26 103
use NAND2X1  _53_
timestamp 1590258663
transform 1 0 396 0 1 105
box -2 -3 26 103
use NOR2X1  _88_
timestamp 1590258663
transform 1 0 420 0 1 105
box -2 -3 26 103
use NAND2X1  _60_
timestamp 1590258663
transform -1 0 468 0 -1 105
box -2 -3 26 103
use NAND2X1  _89_
timestamp 1590258663
transform 1 0 444 0 1 105
box -2 -3 26 103
use FILL  SFILL4680x50
timestamp 1590258663
transform -1 0 476 0 -1 105
box -2 -3 10 103
use FILL  SFILL4760x50
timestamp 1590258663
transform -1 0 484 0 -1 105
box -2 -3 10 103
use FILL  SFILL4840x50
timestamp 1590258663
transform -1 0 492 0 -1 105
box -2 -3 10 103
use FILL  SFILL4680x1050
timestamp 1590258663
transform 1 0 468 0 1 105
box -2 -3 10 103
use FILL  SFILL4760x1050
timestamp 1590258663
transform 1 0 476 0 1 105
box -2 -3 10 103
use FILL  SFILL4840x1050
timestamp 1590258663
transform 1 0 484 0 1 105
box -2 -3 10 103
use NOR2X1  _83_
timestamp 1590258663
transform 1 0 492 0 -1 105
box -2 -3 26 103
use NAND2X1  _84_
timestamp 1590258663
transform -1 0 540 0 -1 105
box -2 -3 26 103
use INVX1  _82_
timestamp 1590258663
transform -1 0 556 0 -1 105
box -2 -3 18 103
use AND2X2  _62_
timestamp 1590258663
transform -1 0 524 0 1 105
box -2 -3 34 103
use INVX1  _49_
timestamp 1590258663
transform 1 0 524 0 1 105
box -2 -3 18 103
use NAND2X1  _51_
timestamp 1590258663
transform 1 0 540 0 1 105
box -2 -3 26 103
use INVX1  _86_
timestamp 1590258663
transform -1 0 572 0 -1 105
box -2 -3 18 103
use XOR2X1  _85_
timestamp 1590258663
transform -1 0 628 0 -1 105
box -2 -3 58 103
use NAND2X1  _50_
timestamp 1590258663
transform -1 0 588 0 1 105
box -2 -3 26 103
use XOR2X1  _31_
timestamp 1590258663
transform 1 0 588 0 1 105
box -2 -3 58 103
use FILL  FILL5800x50
timestamp 1590258663
transform -1 0 636 0 -1 105
box -2 -3 10 103
use FILL  FILL5880x50
timestamp 1590258663
transform -1 0 644 0 -1 105
box -2 -3 10 103
use INVX1  _71_
timestamp 1590258663
transform 1 0 4 0 -1 305
box -2 -3 18 103
use XOR2X1  _70_
timestamp 1590258663
transform 1 0 20 0 -1 305
box -2 -3 58 103
use INVX1  _67_
timestamp 1590258663
transform 1 0 76 0 -1 305
box -2 -3 18 103
use NOR2X1  _68_
timestamp 1590258663
transform -1 0 116 0 -1 305
box -2 -3 26 103
use INVX1  _40_
timestamp 1590258663
transform 1 0 116 0 -1 305
box -2 -3 18 103
use NAND2X1  _69_
timestamp 1590258663
transform 1 0 132 0 -1 305
box -2 -3 26 103
use NAND2X1  _41_
timestamp 1590258663
transform -1 0 180 0 -1 305
box -2 -3 26 103
use FILL  SFILL1800x2050
timestamp 1590258663
transform -1 0 188 0 -1 305
box -2 -3 10 103
use XOR2X1  _28_
timestamp 1590258663
transform -1 0 260 0 -1 305
box -2 -3 58 103
use FILL  SFILL1880x2050
timestamp 1590258663
transform -1 0 196 0 -1 305
box -2 -3 10 103
use FILL  SFILL1960x2050
timestamp 1590258663
transform -1 0 204 0 -1 305
box -2 -3 10 103
use BUFX2  _34_
timestamp 1590258663
transform 1 0 260 0 -1 305
box -2 -3 26 103
use NOR2X1  _64_
timestamp 1590258663
transform -1 0 308 0 -1 305
box -2 -3 26 103
use INVX1  _63_
timestamp 1590258663
transform -1 0 324 0 -1 305
box -2 -3 18 103
use INVX1  _66_
timestamp 1590258663
transform -1 0 340 0 -1 305
box -2 -3 18 103
use XOR2X1  _65_
timestamp 1590258663
transform -1 0 396 0 -1 305
box -2 -3 58 103
use BUFX2  _33_
timestamp 1590258663
transform 1 0 396 0 -1 305
box -2 -3 26 103
use INVX1  _91_
timestamp 1590258663
transform 1 0 420 0 -1 305
box -2 -3 18 103
use XOR2X1  _90_
timestamp 1590258663
transform 1 0 436 0 -1 305
box -2 -3 58 103
use INVX1  _87_
timestamp 1590258663
transform -1 0 532 0 -1 305
box -2 -3 18 103
use XOR2X1  _32_
timestamp 1590258663
transform -1 0 588 0 -1 305
box -2 -3 58 103
use FILL  SFILL4920x2050
timestamp 1590258663
transform -1 0 500 0 -1 305
box -2 -3 10 103
use FILL  SFILL5000x2050
timestamp 1590258663
transform -1 0 508 0 -1 305
box -2 -3 10 103
use FILL  SFILL5080x2050
timestamp 1590258663
transform -1 0 516 0 -1 305
box -2 -3 10 103
use BUFX2  _38_
timestamp 1590258663
transform 1 0 588 0 -1 305
box -2 -3 26 103
use BUFX2  _37_
timestamp 1590258663
transform 1 0 612 0 -1 305
box -2 -3 26 103
use FILL  FILL5880x2050
timestamp 1590258663
transform -1 0 644 0 -1 305
box -2 -3 10 103
<< labels >>
flabel metal6 s 460 -6 484 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal6 s 164 -6 188 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 598 338 602 342 3 FreeSans 24 90 0 0 S[5]
port 2 nsew
flabel metal3 s 670 248 674 252 3 FreeSans 24 90 0 0 S[4]
port 3 nsew
flabel metal2 s 254 338 258 342 3 FreeSans 24 90 0 0 S[3]
port 4 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 S[2]
port 5 nsew
flabel metal2 s 270 338 274 342 3 FreeSans 24 90 0 0 S[1]
port 6 nsew
flabel metal2 s 406 338 410 342 3 FreeSans 24 90 0 0 S[0]
port 7 nsew
flabel metal2 s 518 338 522 342 3 FreeSans 24 90 0 0 X[5]
port 8 nsew
flabel metal2 s 574 -22 578 -18 3 FreeSans 24 270 0 0 X[4]
port 9 nsew
flabel metal2 s 198 -22 202 -18 7 FreeSans 24 270 0 0 X[3]
port 10 nsew
flabel metal3 s -26 138 -22 142 7 FreeSans 24 0 0 0 X[2]
port 11 nsew
flabel metal2 s 78 338 82 342 3 FreeSans 24 90 0 0 X[1]
port 12 nsew
flabel metal2 s 318 338 322 342 3 FreeSans 24 90 0 0 X[0]
port 13 nsew
flabel metal2 s 438 338 442 342 3 FreeSans 24 90 0 0 Y[5]
port 14 nsew
flabel metal3 s 670 48 674 52 3 FreeSans 24 270 0 0 Y[4]
port 15 nsew
flabel metal2 s 214 -22 218 -18 7 FreeSans 24 270 0 0 Y[3]
port 16 nsew
flabel metal3 s -26 158 -22 162 7 FreeSans 24 0 0 0 Y[2]
port 17 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 90 0 0 Y[1]
port 18 nsew
flabel metal2 s 342 338 346 342 3 FreeSans 24 90 0 0 Y[0]
port 19 nsew
flabel metal2 s 350 -22 354 -18 7 FreeSans 24 270 0 0 cout
port 20 nsew
<< end >>
