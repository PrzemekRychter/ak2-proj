VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO adder
   CLASS BLOCK ;
   FOREIGN adder ;
   ORIGIN 2.6000 2.2000 ;
   SIZE 70.0000 BY 36.4000 ;
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 30.2000 64.6000 30.8000 ;
	    RECT 0.6000 28.9000 1.0000 30.2000 ;
	    RECT 3.1000 29.9000 3.5000 30.2000 ;
	    RECT 3.0000 28.2000 3.5000 29.9000 ;
	    RECT 6.1000 28.2000 6.6000 30.2000 ;
	    RECT 7.8000 28.9000 8.2000 30.2000 ;
	    RECT 9.4000 28.9000 9.8000 30.2000 ;
	    RECT 11.0000 28.9000 11.4000 30.2000 ;
	    RECT 11.8000 28.9000 12.2000 30.2000 ;
	    RECT 13.4000 27.9000 13.8000 30.2000 ;
	    RECT 17.4000 27.9000 17.8000 30.2000 ;
	    RECT 21.4000 28.2000 21.9000 30.2000 ;
	    RECT 24.5000 29.9000 24.9000 30.2000 ;
	    RECT 24.5000 28.2000 25.0000 29.9000 ;
	    RECT 27.0000 27.9000 27.4000 30.2000 ;
	    RECT 28.6000 28.9000 29.0000 30.2000 ;
	    RECT 30.2000 28.9000 30.6000 30.2000 ;
	    RECT 31.8000 28.9000 32.2000 30.2000 ;
	    RECT 33.4000 28.9000 33.8000 30.2000 ;
	    RECT 35.0000 28.2000 35.5000 30.2000 ;
	    RECT 38.1000 29.9000 38.5000 30.2000 ;
	    RECT 38.1000 28.2000 38.6000 29.9000 ;
	    RECT 40.6000 27.9000 41.0000 30.2000 ;
	    RECT 42.2000 28.9000 42.6000 30.2000 ;
	    RECT 44.7000 29.9000 45.1000 30.2000 ;
	    RECT 44.6000 28.2000 45.1000 29.9000 ;
	    RECT 47.7000 28.2000 48.2000 30.2000 ;
	    RECT 52.6000 28.9000 53.0000 30.2000 ;
	    RECT 54.2000 28.2000 54.7000 30.2000 ;
	    RECT 57.3000 29.9000 57.7000 30.2000 ;
	    RECT 57.3000 28.2000 57.8000 29.9000 ;
	    RECT 59.8000 27.9000 60.2000 30.2000 ;
	    RECT 62.2000 27.9000 62.6000 30.2000 ;
	    RECT 1.4000 10.8000 1.9000 12.8000 ;
	    RECT 4.5000 11.1000 5.0000 12.8000 ;
	    RECT 4.5000 10.8000 4.9000 11.1000 ;
	    RECT 6.2000 10.8000 6.6000 12.1000 ;
	    RECT 7.8000 10.8000 8.2000 12.1000 ;
	    RECT 9.4000 10.8000 9.8000 13.1000 ;
	    RECT 11.8000 10.8000 12.2000 12.1000 ;
	    RECT 13.4000 10.8000 13.8000 12.1000 ;
	    RECT 14.2000 10.8000 14.6000 13.1000 ;
	    RECT 19.8000 11.1000 20.3000 12.8000 ;
	    RECT 19.9000 10.8000 20.3000 11.1000 ;
	    RECT 22.9000 10.8000 23.4000 12.8000 ;
	    RECT 25.4000 10.8000 25.8000 13.1000 ;
	    RECT 27.0000 10.8000 27.4000 13.1000 ;
	    RECT 29.4000 10.8000 29.8000 13.1000 ;
	    RECT 32.6000 10.8000 33.0000 12.1000 ;
	    RECT 33.4000 10.8000 33.8000 13.1000 ;
	    RECT 35.8000 10.8000 36.2000 12.1000 ;
	    RECT 37.4000 10.8000 37.8000 13.1000 ;
	    RECT 39.8000 10.8000 40.2000 13.1000 ;
	    RECT 42.2000 10.8000 42.6000 12.1000 ;
	    RECT 43.8000 10.8000 44.2000 12.1000 ;
	    RECT 44.6000 10.8000 45.0000 13.1000 ;
	    RECT 50.5000 10.8000 50.9000 13.0000 ;
	    RECT 52.6000 10.8000 53.0000 12.1000 ;
	    RECT 54.2000 10.8000 54.6000 13.1000 ;
	    RECT 58.2000 10.8000 58.6000 13.1000 ;
	    RECT 59.8000 11.1000 60.3000 12.8000 ;
	    RECT 59.9000 10.8000 60.3000 11.1000 ;
	    RECT 62.9000 10.8000 63.4000 12.8000 ;
	    RECT 0.2000 10.2000 64.6000 10.8000 ;
	    RECT 1.4000 7.9000 1.8000 10.2000 ;
	    RECT 3.8000 8.2000 4.3000 10.2000 ;
	    RECT 6.9000 9.9000 7.3000 10.2000 ;
	    RECT 6.9000 8.2000 7.4000 9.9000 ;
	    RECT 8.6000 7.9000 9.0000 10.2000 ;
	    RECT 12.6000 7.9000 13.0000 10.2000 ;
	    RECT 14.2000 8.9000 14.6000 10.2000 ;
	    RECT 18.2000 8.2000 18.7000 10.2000 ;
	    RECT 21.3000 9.9000 21.7000 10.2000 ;
	    RECT 21.3000 8.2000 21.8000 9.9000 ;
	    RECT 23.0000 8.9000 23.4000 10.2000 ;
	    RECT 24.6000 8.9000 25.0000 10.2000 ;
	    RECT 27.5000 8.0000 27.9000 10.2000 ;
	    RECT 29.4000 7.9000 29.8000 10.2000 ;
	    RECT 31.8000 8.9000 32.2000 10.2000 ;
	    RECT 33.4000 8.9000 33.8000 10.2000 ;
	    RECT 35.0000 7.9000 35.4000 10.2000 ;
	    RECT 38.2000 7.9000 38.6000 10.2000 ;
	    RECT 39.8000 8.9000 40.2000 10.2000 ;
	    RECT 42.2000 7.9000 42.6000 10.2000 ;
	    RECT 43.8000 8.9000 44.2000 10.2000 ;
	    RECT 46.2000 7.9000 46.6000 10.2000 ;
	    RECT 49.4000 8.9000 49.8000 10.2000 ;
	    RECT 51.0000 8.9000 51.4000 10.2000 ;
	    RECT 53.4000 7.9000 53.8000 10.2000 ;
	    RECT 55.0000 8.9000 55.4000 10.2000 ;
	    RECT 56.6000 8.9000 57.0000 10.2000 ;
	    RECT 58.2000 8.2000 58.7000 10.2000 ;
	    RECT 61.3000 9.9000 61.7000 10.2000 ;
	    RECT 61.3000 8.2000 61.8000 9.9000 ;
         LAYER metal2 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal3 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal4 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.9000 30.2000 47.5000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.9000 10.2000 47.5000 10.3000 ;
         LAYER metal5 ;
	    RECT 46.9000 30.7000 47.5000 30.8000 ;
	    RECT 46.0000 30.3000 48.4000 30.7000 ;
	    RECT 46.6000 30.2000 47.8000 30.3000 ;
	    RECT 46.9000 10.7000 47.5000 10.8000 ;
	    RECT 46.0000 10.3000 48.4000 10.7000 ;
	    RECT 46.6000 10.2000 47.8000 10.3000 ;
         LAYER metal6 ;
	    RECT 46.0000 -0.6000 48.4000 30.7000 ;
      END
   END gnd
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.6000 20.8000 1.0000 23.1000 ;
	    RECT 3.0000 21.1000 3.5000 24.4000 ;
	    RECT 3.1000 20.8000 3.5000 21.1000 ;
	    RECT 6.1000 20.8000 6.6000 24.4000 ;
	    RECT 7.8000 20.8000 8.2000 23.1000 ;
	    RECT 11.0000 20.8000 11.4000 25.1000 ;
	    RECT 11.8000 20.8000 12.2000 23.1000 ;
	    RECT 13.4000 20.8000 13.8000 23.1000 ;
	    RECT 15.0000 20.8000 15.4000 23.1000 ;
	    RECT 15.8000 20.8000 16.2000 23.1000 ;
	    RECT 17.4000 20.8000 17.8000 23.1000 ;
	    RECT 21.4000 20.8000 21.9000 24.4000 ;
	    RECT 24.5000 21.1000 25.0000 24.4000 ;
	    RECT 24.5000 20.8000 24.9000 21.1000 ;
	    RECT 27.0000 20.8000 27.4000 24.5000 ;
	    RECT 30.2000 20.8000 30.6000 25.1000 ;
	    RECT 31.8000 20.8000 32.2000 23.1000 ;
	    RECT 33.4000 20.8000 33.8000 23.1000 ;
	    RECT 35.0000 20.8000 35.5000 24.4000 ;
	    RECT 38.1000 21.1000 38.6000 24.4000 ;
	    RECT 38.1000 20.8000 38.5000 21.1000 ;
	    RECT 40.6000 20.8000 41.0000 24.5000 ;
	    RECT 42.2000 20.8000 42.6000 23.1000 ;
	    RECT 44.6000 21.1000 45.1000 24.4000 ;
	    RECT 44.7000 20.8000 45.1000 21.1000 ;
	    RECT 47.7000 20.8000 48.2000 24.4000 ;
	    RECT 52.6000 20.8000 53.0000 23.1000 ;
	    RECT 54.2000 20.8000 54.7000 24.4000 ;
	    RECT 57.3000 21.1000 57.8000 24.4000 ;
	    RECT 57.3000 20.8000 57.7000 21.1000 ;
	    RECT 59.8000 20.8000 60.2000 24.5000 ;
	    RECT 62.2000 20.8000 62.6000 24.5000 ;
	    RECT 0.2000 20.2000 64.6000 20.8000 ;
	    RECT 1.4000 16.6000 1.9000 20.2000 ;
	    RECT 4.5000 19.9000 4.9000 20.2000 ;
	    RECT 4.5000 16.6000 5.0000 19.9000 ;
	    RECT 6.2000 17.9000 6.6000 20.2000 ;
	    RECT 7.8000 17.9000 8.2000 20.2000 ;
	    RECT 9.4000 17.9000 9.8000 20.2000 ;
	    RECT 11.0000 17.9000 11.4000 20.2000 ;
	    RECT 11.8000 15.9000 12.2000 20.2000 ;
	    RECT 14.2000 17.9000 14.6000 20.2000 ;
	    RECT 15.8000 17.9000 16.2000 20.2000 ;
	    RECT 19.9000 19.9000 20.3000 20.2000 ;
	    RECT 19.8000 16.6000 20.3000 19.9000 ;
	    RECT 22.9000 16.6000 23.4000 20.2000 ;
	    RECT 25.4000 16.5000 25.8000 20.2000 ;
	    RECT 27.0000 17.9000 27.4000 20.2000 ;
	    RECT 28.6000 17.9000 29.0000 20.2000 ;
	    RECT 29.4000 17.9000 29.8000 20.2000 ;
	    RECT 31.0000 17.9000 31.4000 20.2000 ;
	    RECT 32.6000 17.9000 33.0000 20.2000 ;
	    RECT 33.4000 17.9000 33.8000 20.2000 ;
	    RECT 35.0000 17.9000 35.4000 20.2000 ;
	    RECT 35.8000 17.9000 36.2000 20.2000 ;
	    RECT 37.4000 17.9000 37.8000 20.2000 ;
	    RECT 39.0000 17.9000 39.4000 20.2000 ;
	    RECT 39.8000 17.9000 40.2000 20.2000 ;
	    RECT 41.4000 17.9000 41.8000 20.2000 ;
	    RECT 42.2000 15.9000 42.6000 20.2000 ;
	    RECT 44.6000 17.9000 45.0000 20.2000 ;
	    RECT 46.2000 17.9000 46.6000 20.2000 ;
	    RECT 50.2000 16.1000 50.6000 20.2000 ;
	    RECT 51.8000 17.9000 52.2000 20.2000 ;
	    RECT 52.6000 17.9000 53.0000 20.2000 ;
	    RECT 54.2000 17.9000 54.6000 20.2000 ;
	    RECT 55.8000 17.9000 56.2000 20.2000 ;
	    RECT 56.6000 17.9000 57.0000 20.2000 ;
	    RECT 58.2000 17.9000 58.6000 20.2000 ;
	    RECT 59.9000 19.9000 60.3000 20.2000 ;
	    RECT 59.8000 16.6000 60.3000 19.9000 ;
	    RECT 62.9000 16.6000 63.4000 20.2000 ;
	    RECT 1.4000 0.8000 1.8000 4.5000 ;
	    RECT 3.8000 0.8000 4.3000 4.4000 ;
	    RECT 6.9000 1.1000 7.4000 4.4000 ;
	    RECT 6.9000 0.8000 7.3000 1.1000 ;
	    RECT 8.6000 0.8000 9.0000 3.1000 ;
	    RECT 10.2000 0.8000 10.6000 3.1000 ;
	    RECT 11.0000 0.8000 11.4000 3.1000 ;
	    RECT 12.6000 0.8000 13.0000 3.1000 ;
	    RECT 14.2000 0.8000 14.6000 3.1000 ;
	    RECT 18.2000 0.8000 18.7000 4.4000 ;
	    RECT 21.3000 1.1000 21.8000 4.4000 ;
	    RECT 21.3000 0.8000 21.7000 1.1000 ;
	    RECT 23.0000 0.8000 23.4000 3.1000 ;
	    RECT 24.6000 0.8000 25.0000 3.1000 ;
	    RECT 26.2000 0.8000 26.6000 3.1000 ;
	    RECT 27.8000 0.8000 28.2000 4.9000 ;
	    RECT 29.4000 0.8000 29.8000 3.1000 ;
	    RECT 31.0000 0.8000 31.4000 3.1000 ;
	    RECT 31.8000 0.8000 32.2000 5.1000 ;
	    RECT 35.0000 0.8000 35.4000 4.5000 ;
	    RECT 36.6000 0.8000 37.0000 3.1000 ;
	    RECT 38.2000 0.8000 38.6000 3.1000 ;
	    RECT 39.8000 0.8000 40.2000 3.1000 ;
	    RECT 40.6000 0.8000 41.0000 3.1000 ;
	    RECT 42.2000 0.8000 42.6000 3.1000 ;
	    RECT 43.8000 0.8000 44.2000 3.1000 ;
	    RECT 44.6000 0.8000 45.0000 3.1000 ;
	    RECT 46.2000 0.8000 46.6000 3.1000 ;
	    RECT 49.4000 0.8000 49.8000 5.1000 ;
	    RECT 51.8000 0.8000 52.2000 3.1000 ;
	    RECT 53.4000 0.8000 53.8000 3.1000 ;
	    RECT 55.0000 0.8000 55.4000 3.1000 ;
	    RECT 56.6000 0.8000 57.0000 3.1000 ;
	    RECT 58.2000 0.8000 58.7000 4.4000 ;
	    RECT 61.3000 1.1000 61.8000 4.4000 ;
	    RECT 61.3000 0.8000 61.7000 1.1000 ;
	    RECT 0.2000 0.2000 64.6000 0.8000 ;
         LAYER metal2 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal3 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal4 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.3000 20.2000 17.9000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.3000 0.2000 17.9000 0.3000 ;
         LAYER metal5 ;
	    RECT 17.3000 20.7000 17.9000 20.8000 ;
	    RECT 16.4000 20.3000 18.8000 20.7000 ;
	    RECT 17.0000 20.2000 18.2000 20.3000 ;
	    RECT 17.3000 0.7000 17.9000 0.8000 ;
	    RECT 16.4000 0.3000 18.8000 0.7000 ;
	    RECT 17.0000 0.2000 18.2000 0.3000 ;
         LAYER metal6 ;
	    RECT 16.4000 -0.6000 18.8000 30.7000 ;
      END
   END vdd
   PIN S[5]
      PORT
         LAYER metal1 ;
	    RECT 60.6000 26.2000 61.0000 29.9000 ;
	    RECT 60.7000 25.1000 61.0000 26.2000 ;
	    RECT 60.6000 21.1000 61.0000 25.1000 ;
         LAYER metal2 ;
	    RECT 59.8000 34.1000 60.2000 34.2000 ;
	    RECT 59.8000 33.8000 60.9000 34.1000 ;
	    RECT 60.6000 29.2000 60.9000 33.8000 ;
	    RECT 60.6000 28.8000 61.0000 29.2000 ;
      END
   END S[5]
   PIN S[4]
      PORT
         LAYER metal1 ;
	    RECT 63.0000 26.2000 63.4000 29.9000 ;
	    RECT 63.1000 25.1000 63.4000 26.2000 ;
	    RECT 63.0000 24.1000 63.4000 25.1000 ;
	    RECT 64.6000 24.1000 65.0000 24.2000 ;
	    RECT 63.0000 23.8000 65.0000 24.1000 ;
	    RECT 63.0000 21.1000 63.4000 23.8000 ;
         LAYER metal2 ;
	    RECT 64.6000 24.8000 65.0000 25.2000 ;
	    RECT 64.6000 24.2000 64.9000 24.8000 ;
	    RECT 64.6000 23.8000 65.0000 24.2000 ;
         LAYER metal3 ;
	    RECT 64.6000 25.1000 65.0000 25.2000 ;
	    RECT 67.0000 25.1000 67.4000 25.2000 ;
	    RECT 64.6000 24.8000 67.4000 25.1000 ;
      END
   END S[4]
   PIN S[3]
      PORT
         LAYER metal1 ;
	    RECT 26.2000 15.9000 26.6000 19.9000 ;
	    RECT 26.3000 14.8000 26.6000 15.9000 ;
	    RECT 26.2000 11.1000 26.6000 14.8000 ;
         LAYER metal2 ;
	    RECT 25.4000 33.8000 25.8000 34.2000 ;
	    RECT 25.4000 31.2000 25.7000 33.8000 ;
	    RECT 25.4000 30.8000 25.8000 31.2000 ;
	    RECT 26.2000 23.8000 26.6000 24.2000 ;
	    RECT 26.2000 19.2000 26.5000 23.8000 ;
	    RECT 26.2000 18.8000 26.6000 19.2000 ;
         LAYER metal3 ;
	    RECT 25.4000 31.1000 25.8000 31.2000 ;
	    RECT 26.2000 31.1000 26.6000 31.2000 ;
	    RECT 25.4000 30.8000 26.6000 31.1000 ;
	    RECT 25.4000 24.1000 25.8000 24.2000 ;
	    RECT 26.2000 24.1000 26.6000 24.2000 ;
	    RECT 25.4000 23.8000 26.6000 24.1000 ;
         LAYER metal4 ;
	    RECT 26.2000 31.1000 26.6000 31.2000 ;
	    RECT 25.4000 30.8000 26.6000 31.1000 ;
	    RECT 25.4000 24.2000 25.7000 30.8000 ;
	    RECT 25.4000 23.8000 25.8000 24.2000 ;
      END
   END S[3]
   PIN S[2]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 6.2000 1.0000 9.9000 ;
	    RECT 0.6000 5.1000 0.9000 6.2000 ;
	    RECT 0.6000 1.1000 1.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 4.8000 1.0000 5.2000 ;
	    RECT 0.6000 4.2000 0.9000 4.8000 ;
	    RECT 0.6000 3.8000 1.0000 4.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 5.1000 -2.2000 5.2000 ;
	    RECT 0.6000 5.1000 1.0000 5.2000 ;
	    RECT -2.6000 4.8000 1.0000 5.1000 ;
      END
   END S[2]
   PIN S[1]
      PORT
         LAYER metal1 ;
	    RECT 27.8000 26.2000 28.2000 29.9000 ;
	    RECT 27.9000 25.1000 28.2000 26.2000 ;
	    RECT 27.8000 21.1000 28.2000 25.1000 ;
         LAYER metal2 ;
	    RECT 27.0000 34.1000 27.4000 34.2000 ;
	    RECT 27.0000 33.8000 28.1000 34.1000 ;
	    RECT 27.8000 29.2000 28.1000 33.8000 ;
	    RECT 27.8000 28.8000 28.2000 29.2000 ;
      END
   END S[1]
   PIN S[0]
      PORT
         LAYER metal1 ;
	    RECT 41.4000 26.2000 41.8000 29.9000 ;
	    RECT 41.5000 25.1000 41.8000 26.2000 ;
	    RECT 41.4000 21.1000 41.8000 25.1000 ;
         LAYER metal2 ;
	    RECT 40.6000 34.1000 41.0000 34.2000 ;
	    RECT 40.6000 33.8000 41.7000 34.1000 ;
	    RECT 41.4000 29.2000 41.7000 33.8000 ;
	    RECT 41.4000 28.8000 41.8000 29.2000 ;
      END
   END S[0]
   PIN X[5]
      PORT
         LAYER metal1 ;
	    RECT 52.6000 27.8000 53.0000 28.6000 ;
	    RECT 48.2000 26.8000 49.0000 27.2000 ;
         LAYER metal2 ;
	    RECT 51.8000 34.1000 52.2000 34.2000 ;
	    RECT 51.8000 33.8000 52.9000 34.1000 ;
	    RECT 52.6000 28.2000 52.9000 33.8000 ;
	    RECT 48.6000 27.8000 49.0000 28.2000 ;
	    RECT 52.6000 27.8000 53.0000 28.2000 ;
	    RECT 48.6000 27.2000 48.9000 27.8000 ;
	    RECT 48.6000 26.8000 49.0000 27.2000 ;
         LAYER metal3 ;
	    RECT 48.6000 28.1000 49.0000 28.2000 ;
	    RECT 52.6000 28.1000 53.0000 28.2000 ;
	    RECT 48.6000 27.8000 53.0000 28.1000 ;
      END
   END X[5]
   PIN X[4]
      PORT
         LAYER metal1 ;
	    RECT 55.0000 7.8000 55.4000 8.6000 ;
	    RECT 57.4000 6.8000 58.2000 7.2000 ;
         LAYER metal2 ;
	    RECT 55.0000 7.8000 55.4000 8.2000 ;
	    RECT 55.0000 7.2000 55.3000 7.8000 ;
	    RECT 55.0000 6.8000 55.4000 7.2000 ;
	    RECT 56.6000 7.1000 57.0000 7.2000 ;
	    RECT 57.4000 7.1000 57.8000 7.2000 ;
	    RECT 56.6000 6.8000 57.8000 7.1000 ;
	    RECT 57.4000 -1.8000 57.7000 6.8000 ;
	    RECT 57.4000 -2.2000 57.8000 -1.8000 ;
         LAYER metal3 ;
	    RECT 55.0000 7.1000 55.4000 7.2000 ;
	    RECT 56.6000 7.1000 57.0000 7.2000 ;
	    RECT 55.0000 6.8000 57.0000 7.1000 ;
      END
   END X[4]
   PIN X[3]
      PORT
         LAYER metal1 ;
	    RECT 23.0000 7.8000 23.4000 8.6000 ;
	    RECT 17.4000 6.8000 18.2000 7.2000 ;
         LAYER metal2 ;
	    RECT 17.4000 7.8000 17.8000 8.2000 ;
	    RECT 23.0000 7.8000 23.4000 8.2000 ;
	    RECT 17.4000 7.2000 17.7000 7.8000 ;
	    RECT 23.0000 7.2000 23.3000 7.8000 ;
	    RECT 17.4000 6.8000 17.8000 7.2000 ;
	    RECT 23.0000 6.8000 23.4000 7.2000 ;
	    RECT 17.4000 2.2000 17.7000 6.8000 ;
	    RECT 17.4000 1.8000 17.8000 2.2000 ;
	    RECT 19.8000 1.8000 20.2000 2.2000 ;
	    RECT 19.8000 -1.8000 20.1000 1.8000 ;
	    RECT 19.8000 -2.2000 20.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 17.4000 7.8000 17.8000 8.2000 ;
	    RECT 17.4000 7.1000 17.7000 7.8000 ;
	    RECT 23.0000 7.1000 23.4000 7.2000 ;
	    RECT 17.4000 6.8000 23.4000 7.1000 ;
	    RECT 17.4000 2.1000 17.8000 2.2000 ;
	    RECT 19.8000 2.1000 20.2000 2.2000 ;
	    RECT 17.4000 1.8000 20.2000 2.1000 ;
      END
   END X[3]
   PIN X[2]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 13.8000 1.4000 14.2000 ;
	    RECT 7.8000 12.4000 8.2000 13.2000 ;
         LAYER metal2 ;
	    RECT 0.6000 14.8000 1.0000 15.2000 ;
	    RECT 0.6000 14.2000 0.9000 14.8000 ;
	    RECT 0.6000 13.8000 1.0000 14.2000 ;
	    RECT 7.8000 13.8000 8.2000 14.2000 ;
	    RECT 7.8000 13.2000 8.1000 13.8000 ;
	    RECT 7.8000 12.8000 8.2000 13.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 14.8000 1.0000 15.2000 ;
	    RECT -2.6000 14.1000 -2.2000 14.2000 ;
	    RECT 0.6000 14.1000 0.9000 14.8000 ;
	    RECT 7.8000 14.1000 8.2000 14.2000 ;
	    RECT -2.6000 13.8000 8.2000 14.1000 ;
      END
   END X[2]
   PIN X[1]
      PORT
         LAYER metal1 ;
	    RECT 7.8000 27.8000 8.2000 28.6000 ;
	    RECT 6.6000 27.1000 7.4000 27.2000 ;
	    RECT 7.8000 27.1000 8.1000 27.8000 ;
	    RECT 6.6000 26.8000 8.1000 27.1000 ;
         LAYER metal2 ;
	    RECT 7.8000 33.8000 8.2000 34.2000 ;
	    RECT 7.8000 28.2000 8.1000 33.8000 ;
	    RECT 7.8000 27.8000 8.2000 28.2000 ;
      END
   END X[1]
   PIN X[0]
      PORT
         LAYER metal1 ;
	    RECT 31.8000 27.8000 32.2000 28.6000 ;
	    RECT 34.2000 26.8000 35.0000 27.2000 ;
         LAYER metal2 ;
	    RECT 31.8000 33.8000 32.2000 34.2000 ;
	    RECT 31.8000 28.2000 32.1000 33.8000 ;
	    RECT 31.8000 27.8000 32.2000 28.2000 ;
	    RECT 31.8000 27.2000 32.1000 27.8000 ;
	    RECT 31.8000 26.8000 32.2000 27.2000 ;
	    RECT 33.4000 27.1000 33.8000 27.2000 ;
	    RECT 34.2000 27.1000 34.6000 27.2000 ;
	    RECT 33.4000 26.8000 34.6000 27.1000 ;
         LAYER metal3 ;
	    RECT 31.8000 27.1000 32.2000 27.2000 ;
	    RECT 33.4000 27.1000 33.8000 27.2000 ;
	    RECT 31.8000 26.8000 33.8000 27.1000 ;
      END
   END X[0]
   PIN Y[5]
      PORT
         LAYER metal1 ;
	    RECT 42.2000 27.8000 42.6000 28.6000 ;
	    RECT 43.8000 27.1000 44.6000 27.2000 ;
	    RECT 43.8000 27.0000 44.9000 27.1000 ;
	    RECT 43.8000 26.8000 46.0000 27.0000 ;
	    RECT 44.6000 26.7000 46.0000 26.8000 ;
	    RECT 45.6000 26.6000 46.0000 26.7000 ;
         LAYER metal2 ;
	    RECT 43.8000 33.8000 44.2000 34.2000 ;
	    RECT 43.8000 28.2000 44.1000 33.8000 ;
	    RECT 42.2000 28.1000 42.6000 28.2000 ;
	    RECT 43.0000 28.1000 43.4000 28.2000 ;
	    RECT 42.2000 27.8000 43.4000 28.1000 ;
	    RECT 43.8000 27.8000 44.2000 28.2000 ;
	    RECT 43.8000 27.2000 44.1000 27.8000 ;
	    RECT 43.8000 26.8000 44.2000 27.2000 ;
         LAYER metal3 ;
	    RECT 43.0000 28.1000 43.4000 28.2000 ;
	    RECT 43.8000 28.1000 44.2000 28.2000 ;
	    RECT 43.0000 27.8000 44.2000 28.1000 ;
      END
   END Y[5]
   PIN Y[4]
      PORT
         LAYER metal1 ;
	    RECT 56.6000 7.8000 57.0000 8.6000 ;
	    RECT 61.8000 7.1000 62.6000 7.2000 ;
	    RECT 64.6000 7.1000 65.0000 7.2000 ;
	    RECT 61.5000 7.0000 65.0000 7.1000 ;
	    RECT 60.4000 6.8000 65.0000 7.0000 ;
	    RECT 60.4000 6.7000 61.8000 6.8000 ;
	    RECT 60.4000 6.6000 60.8000 6.7000 ;
         LAYER metal2 ;
	    RECT 55.8000 8.1000 56.2000 8.2000 ;
	    RECT 56.6000 8.1000 57.0000 8.2000 ;
	    RECT 55.8000 7.8000 57.0000 8.1000 ;
	    RECT 64.6000 7.8000 65.0000 8.2000 ;
	    RECT 64.6000 7.2000 64.9000 7.8000 ;
	    RECT 64.6000 6.8000 65.0000 7.2000 ;
	    RECT 64.6000 5.2000 64.9000 6.8000 ;
	    RECT 64.6000 4.8000 65.0000 5.2000 ;
         LAYER metal3 ;
	    RECT 55.8000 8.1000 56.2000 8.2000 ;
	    RECT 64.6000 8.1000 65.0000 8.2000 ;
	    RECT 55.8000 7.8000 65.0000 8.1000 ;
	    RECT 64.6000 5.1000 65.0000 5.2000 ;
	    RECT 67.0000 5.1000 67.4000 5.2000 ;
	    RECT 64.6000 4.8000 67.4000 5.1000 ;
      END
   END Y[4]
   PIN Y[3]
      PORT
         LAYER metal1 ;
	    RECT 24.6000 7.8000 25.0000 8.6000 ;
	    RECT 21.8000 7.1000 22.6000 7.2000 ;
	    RECT 21.5000 7.0000 22.6000 7.1000 ;
	    RECT 20.4000 6.8000 22.6000 7.0000 ;
	    RECT 20.4000 6.7000 21.8000 6.8000 ;
	    RECT 20.4000 6.6000 20.8000 6.7000 ;
         LAYER metal2 ;
	    RECT 22.2000 7.8000 22.6000 8.2000 ;
	    RECT 23.8000 8.1000 24.2000 8.2000 ;
	    RECT 24.6000 8.1000 25.0000 8.2000 ;
	    RECT 23.8000 7.8000 25.0000 8.1000 ;
	    RECT 22.2000 7.2000 22.5000 7.8000 ;
	    RECT 22.2000 6.8000 22.6000 7.2000 ;
	    RECT 21.4000 -1.9000 21.8000 -1.8000 ;
	    RECT 22.2000 -1.9000 22.5000 6.8000 ;
	    RECT 21.4000 -2.2000 22.5000 -1.9000 ;
         LAYER metal3 ;
	    RECT 22.2000 8.1000 22.6000 8.2000 ;
	    RECT 23.8000 8.1000 24.2000 8.2000 ;
	    RECT 22.2000 7.8000 24.2000 8.1000 ;
      END
   END Y[3]
   PIN Y[2]
      PORT
         LAYER metal1 ;
	    RECT 3.6000 14.3000 4.0000 14.4000 ;
	    RECT 3.6000 14.2000 5.0000 14.3000 ;
	    RECT 3.6000 14.1000 5.8000 14.2000 ;
	    RECT 3.6000 14.0000 6.5000 14.1000 ;
	    RECT 4.7000 13.9000 6.5000 14.0000 ;
	    RECT 5.0000 13.8000 6.5000 13.9000 ;
	    RECT 6.2000 13.2000 6.5000 13.8000 ;
	    RECT 6.2000 12.4000 6.6000 13.2000 ;
         LAYER metal2 ;
	    RECT 5.4000 15.8000 5.8000 16.2000 ;
	    RECT 5.4000 14.2000 5.7000 15.8000 ;
	    RECT 5.4000 13.8000 5.8000 14.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 16.1000 -2.2000 16.2000 ;
	    RECT 5.4000 16.1000 5.8000 16.2000 ;
	    RECT -2.6000 15.8000 5.8000 16.1000 ;
      END
   END Y[2]
   PIN Y[1]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 27.8000 1.0000 28.6000 ;
	    RECT 2.2000 27.1000 3.0000 27.2000 ;
	    RECT 2.2000 27.0000 3.3000 27.1000 ;
	    RECT 2.2000 26.8000 4.4000 27.0000 ;
	    RECT 3.0000 26.7000 4.4000 26.8000 ;
	    RECT 4.0000 26.6000 4.4000 26.7000 ;
         LAYER metal2 ;
	    RECT 0.6000 27.8000 1.0000 28.2000 ;
	    RECT 0.6000 25.2000 0.9000 27.8000 ;
	    RECT 2.2000 26.8000 2.6000 27.2000 ;
	    RECT 2.2000 25.2000 2.5000 26.8000 ;
	    RECT 0.6000 24.8000 1.0000 25.2000 ;
	    RECT 2.2000 24.8000 2.6000 25.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 25.1000 -2.2000 25.2000 ;
	    RECT 0.6000 25.1000 1.0000 25.2000 ;
	    RECT 2.2000 25.1000 2.6000 25.2000 ;
	    RECT -2.6000 24.8000 2.6000 25.1000 ;
      END
   END Y[1]
   PIN Y[0]
      PORT
         LAYER metal1 ;
	    RECT 33.4000 27.8000 33.8000 28.6000 ;
	    RECT 38.6000 27.1000 39.4000 27.2000 ;
	    RECT 38.3000 27.0000 39.4000 27.1000 ;
	    RECT 37.2000 26.8000 39.4000 27.0000 ;
	    RECT 37.2000 26.7000 38.6000 26.8000 ;
	    RECT 37.2000 26.6000 37.6000 26.7000 ;
         LAYER metal2 ;
	    RECT 34.2000 33.8000 34.6000 34.2000 ;
	    RECT 34.2000 31.2000 34.5000 33.8000 ;
	    RECT 34.2000 31.1000 34.6000 31.2000 ;
	    RECT 33.4000 30.8000 34.6000 31.1000 ;
	    RECT 39.0000 30.8000 39.4000 31.2000 ;
	    RECT 33.4000 28.2000 33.7000 30.8000 ;
	    RECT 33.4000 27.8000 33.8000 28.2000 ;
	    RECT 39.0000 27.2000 39.3000 30.8000 ;
	    RECT 39.0000 26.8000 39.4000 27.2000 ;
         LAYER metal3 ;
	    RECT 34.2000 31.1000 34.6000 31.2000 ;
	    RECT 39.0000 31.1000 39.4000 31.2000 ;
	    RECT 34.2000 30.8000 39.4000 31.1000 ;
      END
   END Y[0]
   PIN cout
      PORT
         LAYER metal1 ;
	    RECT 34.2000 6.2000 34.6000 9.9000 ;
	    RECT 34.2000 5.1000 34.5000 6.2000 ;
	    RECT 34.2000 1.1000 34.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 34.2000 1.8000 34.6000 2.2000 ;
	    RECT 34.2000 -1.9000 34.5000 1.8000 ;
	    RECT 35.0000 -1.9000 35.4000 -1.8000 ;
	    RECT 34.2000 -2.2000 35.4000 -1.9000 ;
      END
   END cout
   OBS
         LAYER metal1 ;
	    RECT 1.4000 21.1000 1.8000 29.9000 ;
	    RECT 2.2000 27.9000 2.6000 29.9000 ;
	    RECT 4.4000 28.1000 5.2000 29.9000 ;
	    RECT 2.2000 27.6000 3.5000 27.9000 ;
	    RECT 3.1000 27.5000 3.5000 27.6000 ;
	    RECT 3.8000 27.4000 4.6000 27.8000 ;
	    RECT 4.9000 27.1000 5.2000 28.1000 ;
	    RECT 7.0000 27.9000 7.4000 29.9000 ;
	    RECT 5.5000 27.4000 5.9000 27.8000 ;
	    RECT 6.2000 27.6000 7.4000 27.9000 ;
	    RECT 6.2000 27.5000 6.6000 27.6000 ;
	    RECT 4.7000 26.8000 5.2000 27.1000 ;
	    RECT 5.6000 27.2000 5.9000 27.4000 ;
	    RECT 5.6000 26.8000 6.0000 27.2000 ;
	    RECT 4.7000 26.2000 5.0000 26.8000 ;
	    RECT 3.3000 26.1000 3.7000 26.2000 ;
	    RECT 3.3000 25.8000 4.1000 26.1000 ;
	    RECT 4.6000 25.8000 5.0000 26.2000 ;
	    RECT 3.7000 25.7000 4.1000 25.8000 ;
	    RECT 4.7000 25.1000 5.0000 25.8000 ;
	    RECT 8.6000 26.1000 9.0000 29.9000 ;
	    RECT 10.2000 28.9000 10.6000 29.9000 ;
	    RECT 10.2000 27.2000 10.5000 28.9000 ;
	    RECT 11.0000 27.8000 11.4000 28.6000 ;
	    RECT 11.8000 27.8000 12.2000 28.6000 ;
	    RECT 10.2000 27.1000 10.6000 27.2000 ;
	    RECT 11.8000 27.1000 12.1000 27.8000 ;
	    RECT 10.2000 26.8000 12.1000 27.1000 ;
	    RECT 9.4000 26.1000 9.8000 26.2000 ;
	    RECT 8.6000 25.8000 9.8000 26.1000 ;
	    RECT 2.2000 24.8000 3.5000 25.1000 ;
	    RECT 2.2000 21.1000 2.6000 24.8000 ;
	    RECT 3.1000 24.7000 3.5000 24.8000 ;
	    RECT 4.4000 21.1000 5.2000 25.1000 ;
	    RECT 6.2000 24.8000 7.4000 25.1000 ;
	    RECT 6.2000 24.7000 6.6000 24.8000 ;
	    RECT 7.0000 21.1000 7.4000 24.8000 ;
	    RECT 8.6000 21.1000 9.0000 25.8000 ;
	    RECT 9.4000 25.4000 9.8000 25.8000 ;
	    RECT 10.2000 25.1000 10.5000 26.8000 ;
	    RECT 9.7000 24.7000 10.6000 25.1000 ;
	    RECT 9.7000 21.1000 10.1000 24.7000 ;
	    RECT 12.6000 21.1000 13.0000 29.9000 ;
	    RECT 14.7000 28.2000 15.1000 29.9000 ;
	    RECT 14.2000 27.9000 15.1000 28.2000 ;
	    RECT 16.1000 28.2000 16.5000 29.9000 ;
	    RECT 16.1000 27.9000 17.0000 28.2000 ;
	    RECT 13.4000 26.8000 13.8000 27.6000 ;
	    RECT 14.2000 26.1000 14.6000 27.9000 ;
	    RECT 14.2000 25.8000 16.1000 26.1000 ;
	    RECT 14.2000 21.1000 14.6000 25.8000 ;
	    RECT 15.8000 25.2000 16.1000 25.8000 ;
	    RECT 15.0000 24.4000 15.4000 25.2000 ;
	    RECT 15.8000 24.4000 16.2000 25.2000 ;
	    RECT 16.6000 21.1000 17.0000 27.9000 ;
	    RECT 20.6000 27.9000 21.0000 29.9000 ;
	    RECT 22.8000 28.1000 23.6000 29.9000 ;
	    RECT 20.6000 27.6000 21.8000 27.9000 ;
	    RECT 17.4000 26.8000 17.8000 27.6000 ;
	    RECT 21.4000 27.5000 21.8000 27.6000 ;
	    RECT 22.1000 27.4000 22.5000 27.8000 ;
	    RECT 22.1000 27.2000 22.4000 27.4000 ;
	    RECT 19.0000 27.1000 19.4000 27.2000 ;
	    RECT 20.6000 27.1000 21.4000 27.2000 ;
	    RECT 19.0000 26.8000 21.4000 27.1000 ;
	    RECT 22.0000 26.8000 22.4000 27.2000 ;
	    RECT 22.8000 27.1000 23.1000 28.1000 ;
	    RECT 25.4000 27.9000 25.8000 29.9000 ;
	    RECT 23.4000 27.4000 24.2000 27.8000 ;
	    RECT 24.5000 27.6000 25.8000 27.9000 ;
	    RECT 26.2000 27.6000 26.6000 29.9000 ;
	    RECT 29.4000 28.9000 29.8000 29.9000 ;
	    RECT 24.5000 27.5000 24.9000 27.6000 ;
	    RECT 26.2000 27.3000 27.3000 27.6000 ;
	    RECT 25.0000 27.1000 25.8000 27.2000 ;
	    RECT 22.8000 26.8000 23.3000 27.1000 ;
	    RECT 24.7000 27.0000 25.8000 27.1000 ;
	    RECT 23.0000 26.2000 23.3000 26.8000 ;
	    RECT 23.6000 26.8000 25.8000 27.0000 ;
	    RECT 23.6000 26.7000 25.0000 26.8000 ;
	    RECT 23.6000 26.6000 24.0000 26.7000 ;
	    RECT 25.4000 26.2000 25.7000 26.8000 ;
	    RECT 23.0000 25.8000 23.4000 26.2000 ;
	    RECT 24.3000 26.1000 24.7000 26.2000 ;
	    RECT 23.9000 25.8000 24.7000 26.1000 ;
	    RECT 25.4000 25.8000 25.8000 26.2000 ;
	    RECT 26.2000 25.8000 26.6000 26.6000 ;
	    RECT 27.0000 25.8000 27.3000 27.3000 ;
	    RECT 29.4000 27.2000 29.7000 28.9000 ;
	    RECT 30.2000 27.8000 30.6000 28.6000 ;
	    RECT 29.4000 26.8000 29.8000 27.2000 ;
	    RECT 30.2000 26.8000 30.6000 27.2000 ;
	    RECT 23.0000 25.2000 23.3000 25.8000 ;
	    RECT 23.9000 25.7000 24.3000 25.8000 ;
	    RECT 27.0000 25.4000 27.6000 25.8000 ;
	    RECT 28.6000 25.4000 29.0000 26.2000 ;
	    RECT 23.0000 25.1000 24.2000 25.2000 ;
	    RECT 27.0000 25.1000 27.3000 25.4000 ;
	    RECT 29.4000 25.1000 29.7000 26.8000 ;
	    RECT 30.2000 26.1000 30.5000 26.8000 ;
	    RECT 31.0000 26.1000 31.4000 29.9000 ;
	    RECT 30.2000 25.8000 31.4000 26.1000 ;
	    RECT 20.6000 24.8000 21.8000 25.1000 ;
	    RECT 20.6000 21.1000 21.0000 24.8000 ;
	    RECT 21.4000 24.7000 21.8000 24.8000 ;
	    RECT 22.8000 24.8000 24.2000 25.1000 ;
	    RECT 24.5000 24.8000 25.8000 25.1000 ;
	    RECT 22.8000 21.1000 23.6000 24.8000 ;
	    RECT 24.5000 24.7000 24.9000 24.8000 ;
	    RECT 25.4000 21.1000 25.8000 24.8000 ;
	    RECT 26.2000 24.8000 27.3000 25.1000 ;
	    RECT 26.2000 21.1000 26.6000 24.8000 ;
	    RECT 28.9000 24.7000 29.8000 25.1000 ;
	    RECT 28.9000 21.1000 29.3000 24.7000 ;
	    RECT 31.0000 21.1000 31.4000 25.8000 ;
	    RECT 32.6000 21.1000 33.0000 29.9000 ;
	    RECT 34.2000 27.9000 34.6000 29.9000 ;
	    RECT 36.4000 28.1000 37.2000 29.9000 ;
	    RECT 34.2000 27.6000 35.4000 27.9000 ;
	    RECT 35.0000 27.5000 35.4000 27.6000 ;
	    RECT 35.7000 27.4000 36.1000 27.8000 ;
	    RECT 35.7000 27.2000 36.0000 27.4000 ;
	    RECT 35.6000 26.8000 36.0000 27.2000 ;
	    RECT 36.4000 27.1000 36.7000 28.1000 ;
	    RECT 39.0000 27.9000 39.4000 29.9000 ;
	    RECT 37.0000 27.4000 37.8000 27.8000 ;
	    RECT 38.1000 27.6000 39.4000 27.9000 ;
	    RECT 39.8000 27.6000 40.2000 29.9000 ;
	    RECT 38.1000 27.5000 38.5000 27.6000 ;
	    RECT 39.8000 27.3000 40.9000 27.6000 ;
	    RECT 36.4000 26.8000 36.9000 27.1000 ;
	    RECT 36.6000 26.2000 36.9000 26.8000 ;
	    RECT 36.6000 25.8000 37.0000 26.2000 ;
	    RECT 37.9000 26.1000 38.3000 26.2000 ;
	    RECT 37.5000 25.8000 38.3000 26.1000 ;
	    RECT 39.0000 26.1000 39.4000 26.2000 ;
	    RECT 39.8000 26.1000 40.2000 26.6000 ;
	    RECT 39.0000 25.8000 40.2000 26.1000 ;
	    RECT 40.6000 25.8000 40.9000 27.3000 ;
	    RECT 36.6000 25.1000 36.9000 25.8000 ;
	    RECT 37.5000 25.7000 37.9000 25.8000 ;
	    RECT 40.6000 25.4000 41.2000 25.8000 ;
	    RECT 40.6000 25.1000 40.9000 25.4000 ;
	    RECT 34.2000 24.8000 35.4000 25.1000 ;
	    RECT 34.2000 21.1000 34.6000 24.8000 ;
	    RECT 35.0000 24.7000 35.4000 24.8000 ;
	    RECT 36.4000 21.1000 37.2000 25.1000 ;
	    RECT 38.1000 24.8000 39.4000 25.1000 ;
	    RECT 38.1000 24.7000 38.5000 24.8000 ;
	    RECT 39.0000 21.1000 39.4000 24.8000 ;
	    RECT 39.8000 24.8000 40.9000 25.1000 ;
	    RECT 39.8000 21.1000 40.2000 24.8000 ;
	    RECT 42.2000 24.1000 42.6000 24.2000 ;
	    RECT 43.0000 24.1000 43.4000 29.9000 ;
	    RECT 43.8000 27.9000 44.2000 29.9000 ;
	    RECT 46.0000 28.1000 46.8000 29.9000 ;
	    RECT 43.8000 27.6000 45.1000 27.9000 ;
	    RECT 44.7000 27.5000 45.1000 27.6000 ;
	    RECT 45.4000 27.4000 46.2000 27.8000 ;
	    RECT 46.5000 27.1000 46.8000 28.1000 ;
	    RECT 48.6000 27.9000 49.0000 29.9000 ;
	    RECT 47.1000 27.4000 47.5000 27.8000 ;
	    RECT 47.8000 27.6000 49.0000 27.9000 ;
	    RECT 47.8000 27.5000 48.2000 27.6000 ;
	    RECT 46.3000 26.8000 46.8000 27.1000 ;
	    RECT 47.2000 27.2000 47.5000 27.4000 ;
	    RECT 47.2000 26.8000 47.6000 27.2000 ;
	    RECT 46.3000 26.2000 46.6000 26.8000 ;
	    RECT 44.9000 26.1000 45.3000 26.2000 ;
	    RECT 44.9000 25.8000 45.7000 26.1000 ;
	    RECT 46.2000 25.8000 46.6000 26.2000 ;
	    RECT 45.3000 25.7000 45.7000 25.8000 ;
	    RECT 46.3000 25.1000 46.6000 25.8000 ;
	    RECT 42.2000 23.8000 43.4000 24.1000 ;
	    RECT 43.0000 21.1000 43.4000 23.8000 ;
	    RECT 43.8000 24.8000 45.1000 25.1000 ;
	    RECT 43.8000 21.1000 44.2000 24.8000 ;
	    RECT 44.7000 24.7000 45.1000 24.8000 ;
	    RECT 46.0000 21.1000 46.8000 25.1000 ;
	    RECT 47.8000 24.8000 49.0000 25.1000 ;
	    RECT 47.8000 24.7000 48.2000 24.8000 ;
	    RECT 48.6000 21.1000 49.0000 24.8000 ;
	    RECT 50.2000 22.1000 50.6000 22.2000 ;
	    RECT 51.8000 22.1000 52.2000 29.9000 ;
	    RECT 53.4000 27.9000 53.8000 29.9000 ;
	    RECT 55.6000 28.1000 56.4000 29.9000 ;
	    RECT 53.4000 27.6000 54.6000 27.9000 ;
	    RECT 54.2000 27.5000 54.6000 27.6000 ;
	    RECT 54.9000 27.4000 55.3000 27.8000 ;
	    RECT 54.9000 27.2000 55.2000 27.4000 ;
	    RECT 52.6000 27.1000 53.0000 27.2000 ;
	    RECT 53.4000 27.1000 54.2000 27.2000 ;
	    RECT 52.6000 26.8000 54.2000 27.1000 ;
	    RECT 54.8000 26.8000 55.2000 27.2000 ;
	    RECT 55.6000 27.1000 55.9000 28.1000 ;
	    RECT 58.2000 27.9000 58.6000 29.9000 ;
	    RECT 56.2000 27.4000 57.0000 27.8000 ;
	    RECT 57.3000 27.6000 58.6000 27.9000 ;
	    RECT 59.0000 27.6000 59.4000 29.9000 ;
	    RECT 61.4000 27.6000 61.8000 29.9000 ;
	    RECT 57.3000 27.5000 57.7000 27.6000 ;
	    RECT 59.0000 27.3000 60.1000 27.6000 ;
	    RECT 61.4000 27.3000 62.5000 27.6000 ;
	    RECT 57.8000 27.1000 58.6000 27.2000 ;
	    RECT 55.6000 26.8000 56.1000 27.1000 ;
	    RECT 57.5000 27.0000 58.6000 27.1000 ;
	    RECT 55.8000 26.2000 56.1000 26.8000 ;
	    RECT 56.4000 26.8000 58.6000 27.0000 ;
	    RECT 56.4000 26.7000 57.8000 26.8000 ;
	    RECT 56.4000 26.6000 56.8000 26.7000 ;
	    RECT 55.8000 25.8000 56.2000 26.2000 ;
	    RECT 57.1000 26.1000 57.5000 26.2000 ;
	    RECT 56.7000 25.8000 57.5000 26.1000 ;
	    RECT 59.0000 25.8000 59.4000 26.6000 ;
	    RECT 59.8000 25.8000 60.1000 27.3000 ;
	    RECT 61.4000 25.8000 61.8000 26.6000 ;
	    RECT 62.2000 25.8000 62.5000 27.3000 ;
	    RECT 55.8000 25.2000 56.1000 25.8000 ;
	    RECT 56.7000 25.7000 57.1000 25.8000 ;
	    RECT 59.8000 25.4000 60.4000 25.8000 ;
	    RECT 62.2000 25.4000 62.8000 25.8000 ;
	    RECT 55.8000 25.1000 57.0000 25.2000 ;
	    RECT 59.8000 25.1000 60.1000 25.4000 ;
	    RECT 62.2000 25.1000 62.5000 25.4000 ;
	    RECT 50.2000 21.8000 52.2000 22.1000 ;
	    RECT 51.8000 21.1000 52.2000 21.8000 ;
	    RECT 53.4000 24.8000 54.6000 25.1000 ;
	    RECT 53.4000 21.1000 53.8000 24.8000 ;
	    RECT 54.2000 24.7000 54.6000 24.8000 ;
	    RECT 55.6000 24.8000 57.0000 25.1000 ;
	    RECT 57.3000 24.8000 58.6000 25.1000 ;
	    RECT 55.6000 21.1000 56.4000 24.8000 ;
	    RECT 57.3000 24.7000 57.7000 24.8000 ;
	    RECT 58.2000 21.1000 58.6000 24.8000 ;
	    RECT 59.0000 24.8000 60.1000 25.1000 ;
	    RECT 61.4000 24.8000 62.5000 25.1000 ;
	    RECT 59.0000 21.1000 59.4000 24.8000 ;
	    RECT 61.4000 21.1000 61.8000 24.8000 ;
	    RECT 0.6000 16.2000 1.0000 19.9000 ;
	    RECT 1.4000 16.2000 1.8000 16.3000 ;
	    RECT 0.6000 15.9000 1.8000 16.2000 ;
	    RECT 2.8000 15.9000 3.6000 19.9000 ;
	    RECT 4.5000 16.2000 4.9000 16.3000 ;
	    RECT 5.4000 16.2000 5.8000 19.9000 ;
	    RECT 4.5000 15.9000 5.8000 16.2000 ;
	    RECT 3.0000 15.2000 3.3000 15.9000 ;
	    RECT 3.9000 15.2000 4.3000 15.3000 ;
	    RECT 3.0000 14.8000 3.4000 15.2000 ;
	    RECT 3.9000 14.9000 4.7000 15.2000 ;
	    RECT 4.3000 14.8000 4.7000 14.9000 ;
	    RECT 3.0000 14.2000 3.3000 14.8000 ;
	    RECT 2.0000 13.8000 2.4000 14.2000 ;
	    RECT 2.1000 13.6000 2.4000 13.8000 ;
	    RECT 2.8000 13.9000 3.3000 14.2000 ;
	    RECT 1.4000 13.4000 1.8000 13.5000 ;
	    RECT 0.6000 13.1000 1.8000 13.4000 ;
	    RECT 2.1000 13.2000 2.5000 13.6000 ;
	    RECT 0.6000 11.1000 1.0000 13.1000 ;
	    RECT 2.8000 12.9000 3.1000 13.9000 ;
	    RECT 3.4000 13.2000 4.2000 13.6000 ;
	    RECT 4.5000 13.4000 4.9000 13.5000 ;
	    RECT 4.5000 13.1000 5.8000 13.4000 ;
	    RECT 2.8000 11.1000 3.6000 12.9000 ;
	    RECT 5.4000 11.1000 5.8000 13.1000 ;
	    RECT 7.0000 11.1000 7.4000 19.9000 ;
	    RECT 8.6000 16.1000 9.0000 19.9000 ;
	    RECT 9.4000 16.8000 9.8000 17.2000 ;
	    RECT 9.4000 16.1000 9.7000 16.8000 ;
	    RECT 8.6000 15.8000 9.7000 16.1000 ;
	    RECT 8.6000 11.1000 9.0000 15.8000 ;
	    RECT 9.4000 13.4000 9.8000 14.2000 ;
	    RECT 10.2000 13.1000 10.6000 19.9000 ;
	    RECT 11.0000 15.8000 11.4000 16.6000 ;
	    RECT 13.1000 16.3000 13.5000 19.9000 ;
	    RECT 12.6000 15.9000 13.5000 16.3000 ;
	    RECT 12.7000 14.2000 13.0000 15.9000 ;
	    RECT 13.4000 14.8000 13.8000 15.6000 ;
	    RECT 12.6000 13.8000 13.0000 14.2000 ;
	    RECT 13.4000 14.1000 13.8000 14.2000 ;
	    RECT 14.2000 14.1000 14.6000 14.2000 ;
	    RECT 13.4000 13.8000 14.6000 14.1000 ;
	    RECT 10.2000 12.8000 11.1000 13.1000 ;
	    RECT 10.7000 11.1000 11.1000 12.8000 ;
	    RECT 11.8000 12.4000 12.2000 13.2000 ;
	    RECT 12.7000 13.1000 13.0000 13.8000 ;
	    RECT 14.2000 13.4000 14.6000 13.8000 ;
	    RECT 13.4000 13.1000 13.8000 13.2000 ;
	    RECT 12.6000 12.8000 13.8000 13.1000 ;
	    RECT 15.0000 13.1000 15.4000 19.9000 ;
	    RECT 15.8000 15.8000 16.2000 16.6000 ;
	    RECT 19.0000 16.2000 19.4000 19.9000 ;
	    RECT 19.9000 16.2000 20.3000 16.3000 ;
	    RECT 19.0000 15.9000 20.3000 16.2000 ;
	    RECT 21.2000 15.9000 22.0000 19.9000 ;
	    RECT 23.0000 16.2000 23.4000 16.3000 ;
	    RECT 23.8000 16.2000 24.2000 19.9000 ;
	    RECT 23.0000 15.9000 24.2000 16.2000 ;
	    RECT 24.6000 16.2000 25.0000 19.9000 ;
	    RECT 24.6000 15.9000 25.7000 16.2000 ;
	    RECT 20.5000 15.2000 20.9000 15.3000 ;
	    RECT 21.5000 15.2000 21.8000 15.9000 ;
	    RECT 25.4000 15.6000 25.7000 15.9000 ;
	    RECT 27.0000 16.1000 27.4000 16.2000 ;
	    RECT 27.8000 16.1000 28.2000 19.9000 ;
	    RECT 29.4000 17.1000 29.8000 17.2000 ;
	    RECT 30.2000 17.1000 30.6000 19.9000 ;
	    RECT 29.4000 16.8000 30.6000 17.1000 ;
	    RECT 27.0000 15.8000 28.2000 16.1000 ;
	    RECT 28.6000 15.8000 29.0000 16.6000 ;
	    RECT 25.4000 15.2000 26.0000 15.6000 ;
	    RECT 20.1000 14.9000 20.9000 15.2000 ;
	    RECT 21.4000 15.1000 21.8000 15.2000 ;
	    RECT 24.6000 15.1000 25.0000 15.2000 ;
	    RECT 20.1000 14.8000 20.5000 14.9000 ;
	    RECT 21.4000 14.8000 25.0000 15.1000 ;
	    RECT 20.8000 14.3000 21.2000 14.4000 ;
	    RECT 19.8000 14.2000 21.2000 14.3000 ;
	    RECT 15.8000 14.1000 16.2000 14.2000 ;
	    RECT 19.0000 14.1000 21.2000 14.2000 ;
	    RECT 15.8000 14.0000 21.2000 14.1000 ;
	    RECT 21.5000 14.2000 21.8000 14.8000 ;
	    RECT 24.6000 14.4000 25.0000 14.8000 ;
	    RECT 15.8000 13.9000 20.1000 14.0000 ;
	    RECT 21.5000 13.9000 22.0000 14.2000 ;
	    RECT 15.8000 13.8000 19.8000 13.9000 ;
	    RECT 19.9000 13.4000 20.3000 13.5000 ;
	    RECT 19.0000 13.1000 20.3000 13.4000 ;
	    RECT 20.6000 13.2000 21.4000 13.6000 ;
	    RECT 15.0000 12.8000 15.9000 13.1000 ;
	    RECT 12.7000 12.1000 13.0000 12.8000 ;
	    RECT 12.6000 11.1000 13.0000 12.1000 ;
	    RECT 15.5000 11.1000 15.9000 12.8000 ;
	    RECT 19.0000 11.1000 19.4000 13.1000 ;
	    RECT 21.7000 12.9000 22.0000 13.9000 ;
	    RECT 22.4000 13.8000 22.8000 14.2000 ;
	    RECT 23.4000 13.8000 24.2000 14.2000 ;
	    RECT 22.4000 13.6000 22.7000 13.8000 ;
	    RECT 25.4000 13.7000 25.7000 15.2000 ;
	    RECT 22.3000 13.2000 22.7000 13.6000 ;
	    RECT 23.0000 13.4000 23.4000 13.5000 ;
	    RECT 24.6000 13.4000 25.7000 13.7000 ;
	    RECT 27.0000 13.4000 27.4000 14.2000 ;
	    RECT 23.0000 13.1000 24.2000 13.4000 ;
	    RECT 21.2000 11.1000 22.0000 12.9000 ;
	    RECT 23.8000 11.1000 24.2000 13.1000 ;
	    RECT 24.6000 11.1000 25.0000 13.4000 ;
	    RECT 27.8000 13.1000 28.2000 15.8000 ;
	    RECT 29.4000 13.4000 29.8000 14.2000 ;
	    RECT 30.2000 13.1000 30.6000 16.8000 ;
	    RECT 31.0000 15.8000 31.4000 16.6000 ;
	    RECT 31.8000 14.1000 32.2000 19.9000 ;
	    RECT 33.4000 14.1000 33.8000 14.2000 ;
	    RECT 31.8000 13.8000 33.8000 14.1000 ;
	    RECT 27.8000 12.8000 28.7000 13.1000 ;
	    RECT 30.2000 12.8000 31.1000 13.1000 ;
	    RECT 28.3000 11.1000 28.7000 12.8000 ;
	    RECT 30.7000 11.1000 31.1000 12.8000 ;
	    RECT 31.8000 11.1000 32.2000 13.8000 ;
	    RECT 33.4000 13.4000 33.8000 13.8000 ;
	    RECT 34.2000 14.1000 34.6000 19.9000 ;
	    RECT 35.0000 15.8000 35.4000 16.6000 ;
	    RECT 36.6000 14.1000 37.0000 19.9000 ;
	    RECT 37.4000 14.1000 37.8000 14.2000 ;
	    RECT 34.2000 13.8000 36.1000 14.1000 ;
	    RECT 32.6000 12.4000 33.0000 13.2000 ;
	    RECT 34.2000 13.1000 34.6000 13.8000 ;
	    RECT 35.8000 13.2000 36.1000 13.8000 ;
	    RECT 36.6000 13.8000 37.8000 14.1000 ;
	    RECT 34.2000 12.8000 35.1000 13.1000 ;
	    RECT 34.7000 11.1000 35.1000 12.8000 ;
	    RECT 35.8000 12.4000 36.2000 13.2000 ;
	    RECT 36.6000 11.1000 37.0000 13.8000 ;
	    RECT 37.4000 13.4000 37.8000 13.8000 ;
	    RECT 38.2000 14.1000 38.6000 19.9000 ;
	    RECT 39.0000 15.8000 39.4000 16.6000 ;
	    RECT 39.8000 14.1000 40.2000 14.2000 ;
	    RECT 38.2000 13.8000 40.2000 14.1000 ;
	    RECT 38.2000 13.1000 38.6000 13.8000 ;
	    RECT 39.8000 13.4000 40.2000 13.8000 ;
	    RECT 40.6000 13.1000 41.0000 19.9000 ;
	    RECT 41.4000 15.8000 41.8000 17.2000 ;
	    RECT 43.5000 16.3000 43.9000 19.9000 ;
	    RECT 43.0000 15.9000 43.9000 16.3000 ;
	    RECT 43.1000 14.2000 43.4000 15.9000 ;
	    RECT 43.8000 14.8000 44.2000 15.6000 ;
	    RECT 43.0000 13.8000 43.4000 14.2000 ;
	    RECT 43.8000 14.1000 44.2000 14.2000 ;
	    RECT 44.6000 14.1000 45.0000 14.2000 ;
	    RECT 43.8000 13.8000 45.0000 14.1000 ;
	    RECT 38.2000 12.8000 39.1000 13.1000 ;
	    RECT 40.6000 12.8000 41.5000 13.1000 ;
	    RECT 38.7000 11.1000 39.1000 12.8000 ;
	    RECT 41.1000 12.2000 41.5000 12.8000 ;
	    RECT 42.2000 12.4000 42.6000 13.2000 ;
	    RECT 43.1000 12.2000 43.4000 13.8000 ;
	    RECT 44.6000 13.4000 45.0000 13.8000 ;
	    RECT 45.4000 13.1000 45.8000 19.9000 ;
	    RECT 46.2000 15.8000 46.6000 16.6000 ;
	    RECT 49.4000 15.9000 49.8000 19.9000 ;
	    RECT 51.0000 17.9000 51.4000 19.9000 ;
	    RECT 49.4000 15.2000 49.7000 15.9000 ;
	    RECT 51.0000 15.8000 51.3000 17.9000 ;
	    RECT 50.1000 15.5000 51.3000 15.8000 ;
	    RECT 49.4000 14.8000 49.8000 15.2000 ;
	    RECT 49.4000 13.1000 49.7000 14.8000 ;
	    RECT 50.1000 13.8000 50.4000 15.5000 ;
	    RECT 51.0000 14.8000 51.4000 15.2000 ;
	    RECT 51.0000 14.4000 51.3000 14.8000 ;
	    RECT 50.8000 14.1000 51.3000 14.4000 ;
	    RECT 50.8000 14.0000 51.2000 14.1000 ;
	    RECT 51.8000 13.8000 52.2000 14.6000 ;
	    RECT 53.4000 14.1000 53.8000 19.9000 ;
	    RECT 54.2000 14.1000 54.6000 14.2000 ;
	    RECT 53.4000 13.8000 54.6000 14.1000 ;
	    RECT 50.0000 13.7000 50.4000 13.8000 ;
	    RECT 50.0000 13.5000 51.5000 13.7000 ;
	    RECT 50.0000 13.4000 52.1000 13.5000 ;
	    RECT 51.2000 13.2000 52.1000 13.4000 ;
	    RECT 51.8000 13.1000 52.1000 13.2000 ;
	    RECT 45.4000 12.8000 46.3000 13.1000 ;
	    RECT 40.6000 11.8000 41.5000 12.2000 ;
	    RECT 41.1000 11.1000 41.5000 11.8000 ;
	    RECT 43.0000 11.1000 43.4000 12.2000 ;
	    RECT 45.9000 11.1000 46.3000 12.8000 ;
	    RECT 49.4000 12.6000 50.1000 13.1000 ;
	    RECT 49.7000 11.1000 50.1000 12.6000 ;
	    RECT 51.8000 11.1000 52.2000 13.1000 ;
	    RECT 52.6000 12.4000 53.0000 13.2000 ;
	    RECT 53.4000 11.1000 53.8000 13.8000 ;
	    RECT 54.2000 13.4000 54.6000 13.8000 ;
	    RECT 55.0000 13.1000 55.4000 19.9000 ;
	    RECT 55.8000 15.8000 56.2000 16.6000 ;
	    RECT 56.6000 15.8000 57.0000 16.6000 ;
	    RECT 55.8000 15.1000 56.1000 15.8000 ;
	    RECT 57.4000 15.1000 57.8000 19.9000 ;
	    RECT 59.0000 16.2000 59.4000 19.9000 ;
	    RECT 59.9000 16.2000 60.3000 16.3000 ;
	    RECT 59.0000 15.9000 60.3000 16.2000 ;
	    RECT 61.2000 15.9000 62.0000 19.9000 ;
	    RECT 63.0000 16.2000 63.4000 16.3000 ;
	    RECT 63.8000 16.2000 64.2000 19.9000 ;
	    RECT 63.0000 15.9000 64.2000 16.2000 ;
	    RECT 60.5000 15.2000 60.9000 15.3000 ;
	    RECT 61.5000 15.2000 61.8000 15.9000 ;
	    RECT 55.8000 14.8000 57.8000 15.1000 ;
	    RECT 57.4000 13.1000 57.8000 14.8000 ;
	    RECT 58.2000 14.8000 58.6000 15.2000 ;
	    RECT 60.1000 14.9000 60.9000 15.2000 ;
	    RECT 60.1000 14.8000 60.5000 14.9000 ;
	    RECT 61.4000 14.8000 61.8000 15.2000 ;
	    RECT 58.2000 14.2000 58.5000 14.8000 ;
	    RECT 60.8000 14.3000 61.2000 14.4000 ;
	    RECT 59.8000 14.2000 61.2000 14.3000 ;
	    RECT 58.2000 14.1000 58.6000 14.2000 ;
	    RECT 59.0000 14.1000 61.2000 14.2000 ;
	    RECT 58.2000 14.0000 61.2000 14.1000 ;
	    RECT 61.5000 14.2000 61.8000 14.8000 ;
	    RECT 58.2000 13.9000 60.1000 14.0000 ;
	    RECT 61.5000 13.9000 62.0000 14.2000 ;
	    RECT 58.2000 13.8000 59.8000 13.9000 ;
	    RECT 58.2000 13.4000 58.6000 13.8000 ;
	    RECT 59.9000 13.4000 60.3000 13.5000 ;
	    RECT 55.0000 12.8000 55.9000 13.1000 ;
	    RECT 55.5000 11.1000 55.9000 12.8000 ;
	    RECT 56.9000 12.8000 57.8000 13.1000 ;
	    RECT 59.0000 13.1000 60.3000 13.4000 ;
	    RECT 60.6000 13.2000 61.4000 13.6000 ;
	    RECT 56.9000 11.1000 57.3000 12.8000 ;
	    RECT 59.0000 11.1000 59.4000 13.1000 ;
	    RECT 61.7000 12.9000 62.0000 13.9000 ;
	    RECT 62.4000 13.8000 62.8000 14.2000 ;
	    RECT 63.4000 13.8000 64.2000 14.2000 ;
	    RECT 62.4000 13.6000 62.7000 13.8000 ;
	    RECT 62.3000 13.2000 62.7000 13.6000 ;
	    RECT 63.0000 13.4000 63.4000 13.5000 ;
	    RECT 63.0000 13.1000 64.2000 13.4000 ;
	    RECT 61.2000 11.1000 62.0000 12.9000 ;
	    RECT 63.8000 11.1000 64.2000 13.1000 ;
	    RECT 2.2000 7.6000 2.6000 9.9000 ;
	    RECT 3.0000 7.9000 3.4000 9.9000 ;
	    RECT 5.2000 8.1000 6.0000 9.9000 ;
	    RECT 3.0000 7.6000 4.2000 7.9000 ;
	    RECT 1.5000 7.3000 2.6000 7.6000 ;
	    RECT 3.8000 7.5000 4.2000 7.6000 ;
	    RECT 4.5000 7.4000 4.9000 7.8000 ;
	    RECT 1.5000 5.8000 1.8000 7.3000 ;
	    RECT 4.5000 7.2000 4.8000 7.4000 ;
	    RECT 3.0000 6.8000 3.8000 7.2000 ;
	    RECT 4.4000 6.8000 4.8000 7.2000 ;
	    RECT 5.2000 7.1000 5.5000 8.1000 ;
	    RECT 7.8000 7.9000 8.2000 9.9000 ;
	    RECT 9.9000 8.2000 10.3000 9.9000 ;
	    RECT 11.3000 9.2000 11.7000 9.9000 ;
	    RECT 11.0000 8.8000 11.7000 9.2000 ;
	    RECT 5.8000 7.4000 6.6000 7.8000 ;
	    RECT 6.9000 7.6000 8.2000 7.9000 ;
	    RECT 9.4000 7.9000 10.3000 8.2000 ;
	    RECT 11.3000 8.2000 11.7000 8.8000 ;
	    RECT 11.3000 7.9000 12.2000 8.2000 ;
	    RECT 6.9000 7.5000 7.3000 7.6000 ;
	    RECT 7.4000 7.1000 8.2000 7.2000 ;
	    RECT 8.6000 7.1000 9.0000 7.6000 ;
	    RECT 5.2000 6.8000 5.7000 7.1000 ;
	    RECT 7.1000 7.0000 9.0000 7.1000 ;
	    RECT 2.2000 6.1000 2.6000 6.6000 ;
	    RECT 5.4000 6.2000 5.7000 6.8000 ;
	    RECT 6.0000 6.8000 9.0000 7.0000 ;
	    RECT 6.0000 6.7000 7.4000 6.8000 ;
	    RECT 6.0000 6.6000 6.4000 6.7000 ;
	    RECT 5.4000 6.1000 5.8000 6.2000 ;
	    RECT 6.7000 6.1000 7.1000 6.2000 ;
	    RECT 2.2000 5.8000 5.8000 6.1000 ;
	    RECT 6.3000 5.8000 7.1000 6.1000 ;
	    RECT 9.4000 6.1000 9.8000 7.9000 ;
	    RECT 9.4000 5.8000 11.3000 6.1000 ;
	    RECT 1.2000 5.4000 1.8000 5.8000 ;
	    RECT 1.5000 5.1000 1.8000 5.4000 ;
	    RECT 5.4000 5.1000 5.7000 5.8000 ;
	    RECT 6.3000 5.7000 6.7000 5.8000 ;
	    RECT 1.5000 4.8000 2.6000 5.1000 ;
	    RECT 2.2000 1.1000 2.6000 4.8000 ;
	    RECT 3.0000 4.8000 4.2000 5.1000 ;
	    RECT 3.0000 1.1000 3.4000 4.8000 ;
	    RECT 3.8000 4.7000 4.2000 4.8000 ;
	    RECT 5.2000 1.1000 6.0000 5.1000 ;
	    RECT 6.9000 4.8000 8.2000 5.1000 ;
	    RECT 6.9000 4.7000 7.3000 4.8000 ;
	    RECT 7.8000 1.1000 8.2000 4.8000 ;
	    RECT 9.4000 1.1000 9.8000 5.8000 ;
	    RECT 11.0000 5.2000 11.3000 5.8000 ;
	    RECT 10.2000 4.4000 10.6000 5.2000 ;
	    RECT 11.0000 4.4000 11.4000 5.2000 ;
	    RECT 11.8000 1.1000 12.2000 7.9000 ;
	    RECT 12.6000 7.1000 13.0000 7.6000 ;
	    RECT 13.4000 7.1000 13.8000 9.9000 ;
	    RECT 14.2000 7.8000 14.6000 8.6000 ;
	    RECT 17.4000 7.9000 17.8000 9.9000 ;
	    RECT 19.6000 8.1000 20.4000 9.9000 ;
	    RECT 17.4000 7.6000 18.6000 7.9000 ;
	    RECT 18.2000 7.5000 18.6000 7.6000 ;
	    RECT 18.9000 7.4000 19.3000 7.8000 ;
	    RECT 18.9000 7.2000 19.2000 7.4000 ;
	    RECT 12.6000 6.8000 13.8000 7.1000 ;
	    RECT 18.8000 6.8000 19.2000 7.2000 ;
	    RECT 19.6000 7.1000 19.9000 8.1000 ;
	    RECT 22.2000 7.9000 22.6000 9.9000 ;
	    RECT 20.2000 7.4000 21.0000 7.8000 ;
	    RECT 21.3000 7.6000 22.6000 7.9000 ;
	    RECT 21.3000 7.5000 21.7000 7.6000 ;
	    RECT 19.6000 6.8000 20.1000 7.1000 ;
	    RECT 13.4000 1.1000 13.8000 6.8000 ;
	    RECT 19.8000 6.2000 20.1000 6.8000 ;
	    RECT 19.8000 5.8000 20.2000 6.2000 ;
	    RECT 21.1000 6.1000 21.5000 6.2000 ;
	    RECT 20.7000 5.8000 21.5000 6.1000 ;
	    RECT 19.8000 5.1000 20.1000 5.8000 ;
	    RECT 20.7000 5.7000 21.1000 5.8000 ;
	    RECT 23.8000 5.1000 24.2000 9.9000 ;
	    RECT 24.6000 5.8000 25.0000 6.2000 ;
	    RECT 24.6000 5.1000 24.9000 5.8000 ;
	    RECT 17.4000 4.8000 18.6000 5.1000 ;
	    RECT 17.4000 1.1000 17.8000 4.8000 ;
	    RECT 18.2000 4.7000 18.6000 4.8000 ;
	    RECT 19.6000 1.1000 20.4000 5.1000 ;
	    RECT 21.3000 4.8000 22.6000 5.1000 ;
	    RECT 21.3000 4.7000 21.7000 4.8000 ;
	    RECT 22.2000 1.1000 22.6000 4.8000 ;
	    RECT 23.8000 4.8000 24.9000 5.1000 ;
	    RECT 23.8000 1.1000 24.2000 4.8000 ;
	    RECT 25.4000 1.1000 25.8000 9.9000 ;
	    RECT 26.2000 7.9000 26.6000 9.9000 ;
	    RECT 28.3000 9.2000 28.7000 9.9000 ;
	    RECT 30.7000 9.2000 31.1000 9.9000 ;
	    RECT 28.3000 8.8000 29.0000 9.2000 ;
	    RECT 30.7000 8.8000 31.4000 9.2000 ;
	    RECT 32.6000 8.8000 33.0000 9.9000 ;
	    RECT 28.3000 8.4000 28.7000 8.8000 ;
	    RECT 28.3000 7.9000 29.0000 8.4000 ;
	    RECT 30.7000 8.2000 31.1000 8.8000 ;
	    RECT 26.3000 7.8000 26.6000 7.9000 ;
	    RECT 26.3000 7.6000 27.2000 7.8000 ;
	    RECT 26.3000 7.5000 28.4000 7.6000 ;
	    RECT 26.9000 7.3000 28.4000 7.5000 ;
	    RECT 28.0000 7.2000 28.4000 7.3000 ;
	    RECT 26.2000 6.4000 26.6000 7.2000 ;
	    RECT 27.2000 6.9000 27.6000 7.0000 ;
	    RECT 27.1000 6.6000 27.6000 6.9000 ;
	    RECT 27.1000 6.2000 27.4000 6.6000 ;
	    RECT 27.0000 5.8000 27.4000 6.2000 ;
	    RECT 28.0000 5.5000 28.3000 7.2000 ;
	    RECT 28.7000 6.2000 29.0000 7.9000 ;
	    RECT 30.2000 7.9000 31.1000 8.2000 ;
	    RECT 29.4000 6.8000 29.8000 7.6000 ;
	    RECT 28.6000 5.8000 29.0000 6.2000 ;
	    RECT 27.1000 5.2000 28.3000 5.5000 ;
	    RECT 27.1000 3.1000 27.4000 5.2000 ;
	    RECT 28.7000 5.1000 29.0000 5.8000 ;
	    RECT 27.0000 1.1000 27.4000 3.1000 ;
	    RECT 28.6000 1.1000 29.0000 5.1000 ;
	    RECT 30.2000 1.1000 30.6000 7.9000 ;
	    RECT 31.8000 7.8000 32.2000 8.6000 ;
	    RECT 32.7000 7.2000 33.0000 8.8000 ;
	    RECT 35.8000 7.6000 36.2000 9.9000 ;
	    RECT 36.9000 8.2000 37.3000 9.9000 ;
	    RECT 36.9000 7.9000 37.8000 8.2000 ;
	    RECT 32.6000 6.8000 33.0000 7.2000 ;
	    RECT 31.0000 4.4000 31.4000 5.2000 ;
	    RECT 32.7000 5.1000 33.0000 6.8000 ;
	    RECT 35.1000 7.3000 36.2000 7.6000 ;
	    RECT 33.4000 5.4000 33.8000 6.2000 ;
	    RECT 35.1000 5.8000 35.4000 7.3000 ;
	    RECT 35.8000 6.1000 36.2000 6.6000 ;
	    RECT 37.4000 6.1000 37.8000 7.9000 ;
	    RECT 38.2000 7.1000 38.6000 7.6000 ;
	    RECT 39.0000 7.1000 39.4000 9.9000 ;
	    RECT 38.2000 6.8000 39.4000 7.1000 ;
	    RECT 39.8000 7.8000 40.2000 8.6000 ;
	    RECT 40.9000 8.2000 41.3000 9.9000 ;
	    RECT 40.9000 7.9000 41.8000 8.2000 ;
	    RECT 39.8000 7.1000 40.1000 7.8000 ;
	    RECT 41.4000 7.1000 41.8000 7.9000 ;
	    RECT 39.8000 6.8000 41.8000 7.1000 ;
	    RECT 42.2000 7.1000 42.6000 7.6000 ;
	    RECT 43.0000 7.1000 43.4000 9.9000 ;
	    RECT 43.8000 7.8000 44.2000 8.6000 ;
	    RECT 44.9000 8.2000 45.3000 9.9000 ;
	    RECT 50.2000 8.9000 50.6000 9.9000 ;
	    RECT 52.1000 9.2000 52.5000 9.9000 ;
	    RECT 44.9000 7.9000 45.8000 8.2000 ;
	    RECT 42.2000 6.8000 43.4000 7.1000 ;
	    RECT 35.8000 5.8000 37.8000 6.1000 ;
	    RECT 34.8000 5.4000 35.4000 5.8000 ;
	    RECT 35.1000 5.1000 35.4000 5.4000 ;
	    RECT 32.6000 4.7000 33.5000 5.1000 ;
	    RECT 35.1000 4.8000 36.2000 5.1000 ;
	    RECT 33.1000 1.1000 33.5000 4.7000 ;
	    RECT 35.8000 1.1000 36.2000 4.8000 ;
	    RECT 36.6000 4.4000 37.0000 5.2000 ;
	    RECT 37.4000 1.1000 37.8000 5.8000 ;
	    RECT 39.0000 1.1000 39.4000 6.8000 ;
	    RECT 40.6000 4.4000 41.0000 5.2000 ;
	    RECT 41.4000 1.1000 41.8000 6.8000 ;
	    RECT 43.0000 1.1000 43.4000 6.8000 ;
	    RECT 44.6000 4.4000 45.0000 5.2000 ;
	    RECT 45.4000 5.1000 45.8000 7.9000 ;
	    RECT 49.4000 7.8000 49.8000 8.6000 ;
	    RECT 46.2000 7.1000 46.6000 7.6000 ;
	    RECT 50.3000 7.2000 50.6000 8.9000 ;
	    RECT 51.8000 8.8000 52.5000 9.2000 ;
	    RECT 52.1000 8.2000 52.5000 8.8000 ;
	    RECT 52.1000 7.9000 53.0000 8.2000 ;
	    RECT 50.2000 7.1000 50.6000 7.2000 ;
	    RECT 51.8000 7.1000 52.2000 7.2000 ;
	    RECT 46.2000 6.8000 52.2000 7.1000 ;
	    RECT 46.2000 5.1000 46.6000 5.2000 ;
	    RECT 50.3000 5.1000 50.6000 6.8000 ;
	    RECT 51.0000 6.1000 51.4000 6.2000 ;
	    RECT 51.0000 5.8000 52.1000 6.1000 ;
	    RECT 51.0000 5.4000 51.4000 5.8000 ;
	    RECT 51.8000 5.2000 52.1000 5.8000 ;
	    RECT 45.4000 4.8000 46.6000 5.1000 ;
	    RECT 45.4000 1.1000 45.8000 4.8000 ;
	    RECT 50.2000 4.7000 51.1000 5.1000 ;
	    RECT 50.7000 1.1000 51.1000 4.7000 ;
	    RECT 51.8000 4.4000 52.2000 5.2000 ;
	    RECT 52.6000 1.1000 53.0000 7.9000 ;
	    RECT 53.4000 6.8000 53.8000 7.6000 ;
	    RECT 54.2000 5.1000 54.6000 9.9000 ;
	    RECT 55.0000 6.1000 55.4000 6.2000 ;
	    RECT 55.8000 6.1000 56.2000 9.9000 ;
	    RECT 57.4000 7.9000 57.8000 9.9000 ;
	    RECT 59.6000 8.1000 60.4000 9.9000 ;
	    RECT 57.4000 7.6000 58.6000 7.9000 ;
	    RECT 58.2000 7.5000 58.6000 7.6000 ;
	    RECT 58.9000 7.4000 59.3000 7.8000 ;
	    RECT 58.9000 7.2000 59.2000 7.4000 ;
	    RECT 58.8000 6.8000 59.2000 7.2000 ;
	    RECT 59.6000 7.1000 59.9000 8.1000 ;
	    RECT 62.2000 7.9000 62.6000 9.9000 ;
	    RECT 60.2000 7.4000 61.0000 7.8000 ;
	    RECT 61.3000 7.6000 62.6000 7.9000 ;
	    RECT 61.3000 7.5000 61.7000 7.6000 ;
	    RECT 59.6000 6.8000 60.1000 7.1000 ;
	    RECT 55.0000 5.8000 56.2000 6.1000 ;
	    RECT 53.4000 4.8000 54.6000 5.1000 ;
	    RECT 53.4000 4.2000 53.7000 4.8000 ;
	    RECT 53.4000 3.8000 53.8000 4.2000 ;
	    RECT 54.2000 1.1000 54.6000 4.8000 ;
	    RECT 55.8000 1.1000 56.2000 5.8000 ;
	    RECT 59.8000 6.2000 60.1000 6.8000 ;
	    RECT 59.8000 5.8000 60.2000 6.2000 ;
	    RECT 61.1000 6.1000 61.5000 6.2000 ;
	    RECT 60.7000 5.8000 61.5000 6.1000 ;
	    RECT 59.8000 5.1000 60.1000 5.8000 ;
	    RECT 60.7000 5.7000 61.1000 5.8000 ;
	    RECT 57.4000 4.8000 58.6000 5.1000 ;
	    RECT 57.4000 1.1000 57.8000 4.8000 ;
	    RECT 58.2000 4.7000 58.6000 4.8000 ;
	    RECT 59.6000 1.1000 60.4000 5.1000 ;
	    RECT 61.3000 4.8000 62.6000 5.1000 ;
	    RECT 61.3000 4.7000 61.7000 4.8000 ;
	    RECT 62.2000 1.1000 62.6000 4.8000 ;
         LAYER metal2 ;
	    RECT 32.6000 28.8000 33.0000 29.2000 ;
	    RECT 32.6000 28.2000 32.9000 28.8000 ;
	    RECT 1.4000 27.8000 1.8000 28.2000 ;
	    RECT 3.1000 27.8000 3.5000 27.9000 ;
	    RECT 1.4000 27.2000 1.7000 27.8000 ;
	    RECT 3.1000 27.5000 5.9000 27.8000 ;
	    RECT 6.2000 27.5000 6.6000 27.9000 ;
	    RECT 1.4000 26.8000 1.8000 27.2000 ;
	    RECT 3.1000 25.1000 3.4000 27.5000 ;
	    RECT 3.8000 27.4000 4.2000 27.5000 ;
	    RECT 5.5000 27.4000 5.9000 27.5000 ;
	    RECT 6.3000 27.1000 6.6000 27.5000 ;
	    RECT 3.8000 26.8000 6.6000 27.1000 ;
	    RECT 11.0000 27.8000 11.4000 28.2000 ;
	    RECT 30.2000 28.1000 30.6000 28.2000 ;
	    RECT 31.0000 28.1000 31.4000 28.2000 ;
	    RECT 11.0000 27.2000 11.3000 27.8000 ;
	    RECT 21.4000 27.5000 21.8000 27.9000 ;
	    RECT 24.5000 27.8000 24.9000 27.9000 ;
	    RECT 30.2000 27.8000 31.4000 28.1000 ;
	    RECT 32.6000 27.8000 33.0000 28.2000 ;
	    RECT 22.1000 27.5000 24.9000 27.8000 ;
	    RECT 11.0000 26.8000 11.4000 27.2000 ;
	    RECT 12.6000 27.1000 13.0000 27.2000 ;
	    RECT 13.4000 27.1000 13.8000 27.2000 ;
	    RECT 12.6000 26.8000 13.8000 27.1000 ;
	    RECT 17.4000 27.1000 17.8000 27.2000 ;
	    RECT 18.2000 27.1000 18.6000 27.2000 ;
	    RECT 17.4000 26.8000 18.6000 27.1000 ;
	    RECT 19.0000 26.8000 19.4000 27.2000 ;
	    RECT 21.4000 27.1000 21.7000 27.5000 ;
	    RECT 22.1000 27.4000 22.5000 27.5000 ;
	    RECT 23.8000 27.4000 24.2000 27.5000 ;
	    RECT 21.4000 26.8000 24.2000 27.1000 ;
	    RECT 3.8000 26.1000 4.1000 26.8000 ;
	    RECT 3.7000 25.7000 4.1000 26.1000 ;
	    RECT 4.6000 26.1000 5.0000 26.2000 ;
	    RECT 5.4000 26.1000 5.8000 26.2000 ;
	    RECT 4.6000 25.8000 5.8000 26.1000 ;
	    RECT 6.3000 25.1000 6.6000 26.8000 ;
	    RECT 19.0000 26.2000 19.3000 26.8000 ;
	    RECT 3.1000 24.7000 3.5000 25.1000 ;
	    RECT 6.2000 24.7000 6.6000 25.1000 ;
	    RECT 9.4000 25.8000 9.8000 26.2000 ;
	    RECT 19.0000 25.8000 19.4000 26.2000 ;
	    RECT 9.4000 25.2000 9.7000 25.8000 ;
	    RECT 9.4000 24.8000 9.8000 25.2000 ;
	    RECT 14.2000 25.1000 14.6000 25.2000 ;
	    RECT 15.0000 25.1000 15.4000 25.2000 ;
	    RECT 14.2000 24.8000 15.4000 25.1000 ;
	    RECT 21.4000 25.1000 21.7000 26.8000 ;
	    RECT 23.9000 26.1000 24.2000 26.8000 ;
	    RECT 23.9000 25.7000 24.3000 26.1000 ;
	    RECT 23.0000 25.1000 23.4000 25.2000 ;
	    RECT 23.8000 25.1000 24.2000 25.2000 ;
	    RECT 24.6000 25.1000 24.9000 27.5000 ;
	    RECT 35.0000 27.5000 35.4000 27.9000 ;
	    RECT 38.1000 27.8000 38.5000 27.9000 ;
	    RECT 35.7000 27.5000 38.5000 27.8000 ;
	    RECT 25.4000 26.8000 25.8000 27.2000 ;
	    RECT 28.6000 27.1000 29.0000 27.2000 ;
	    RECT 29.4000 27.1000 29.8000 27.2000 ;
	    RECT 28.6000 26.8000 29.8000 27.1000 ;
	    RECT 30.2000 26.8000 30.6000 27.2000 ;
	    RECT 35.0000 27.1000 35.3000 27.5000 ;
	    RECT 35.7000 27.4000 36.1000 27.5000 ;
	    RECT 37.4000 27.4000 37.8000 27.5000 ;
	    RECT 35.0000 26.8000 37.8000 27.1000 ;
	    RECT 25.4000 26.2000 25.7000 26.8000 ;
	    RECT 30.2000 26.2000 30.5000 26.8000 ;
	    RECT 25.4000 25.8000 25.8000 26.2000 ;
	    RECT 26.2000 25.8000 26.6000 26.2000 ;
	    RECT 28.6000 26.1000 29.0000 26.2000 ;
	    RECT 29.4000 26.1000 29.8000 26.2000 ;
	    RECT 28.6000 25.8000 29.8000 26.1000 ;
	    RECT 30.2000 25.8000 30.6000 26.2000 ;
	    RECT 21.4000 24.7000 21.8000 25.1000 ;
	    RECT 23.0000 24.8000 24.2000 25.1000 ;
	    RECT 24.5000 24.7000 24.9000 25.1000 ;
	    RECT 26.2000 25.2000 26.5000 25.8000 ;
	    RECT 26.2000 24.8000 26.6000 25.2000 ;
	    RECT 35.0000 25.1000 35.3000 26.8000 ;
	    RECT 35.8000 26.1000 36.2000 26.2000 ;
	    RECT 36.6000 26.1000 37.0000 26.2000 ;
	    RECT 35.8000 25.8000 37.0000 26.1000 ;
	    RECT 37.5000 26.1000 37.8000 26.8000 ;
	    RECT 37.5000 25.7000 37.9000 26.1000 ;
	    RECT 38.2000 25.1000 38.5000 27.5000 ;
	    RECT 44.7000 27.8000 45.1000 27.9000 ;
	    RECT 44.7000 27.5000 47.5000 27.8000 ;
	    RECT 47.8000 27.5000 48.2000 27.9000 ;
	    RECT 39.0000 26.1000 39.4000 26.2000 ;
	    RECT 39.8000 26.1000 40.2000 26.2000 ;
	    RECT 39.0000 25.8000 40.2000 26.1000 ;
	    RECT 35.0000 24.7000 35.4000 25.1000 ;
	    RECT 38.1000 24.7000 38.5000 25.1000 ;
	    RECT 44.7000 25.1000 45.0000 27.5000 ;
	    RECT 45.4000 27.4000 45.8000 27.5000 ;
	    RECT 47.1000 27.4000 47.5000 27.5000 ;
	    RECT 47.9000 27.1000 48.2000 27.5000 ;
	    RECT 54.2000 27.5000 54.6000 27.9000 ;
	    RECT 57.3000 27.8000 57.7000 27.9000 ;
	    RECT 54.9000 27.5000 57.7000 27.8000 ;
	    RECT 45.4000 26.8000 48.2000 27.1000 ;
	    RECT 45.4000 26.1000 45.7000 26.8000 ;
	    RECT 45.3000 25.7000 45.7000 26.1000 ;
	    RECT 46.2000 26.1000 46.6000 26.2000 ;
	    RECT 47.0000 26.1000 47.4000 26.2000 ;
	    RECT 46.2000 25.8000 47.4000 26.1000 ;
	    RECT 47.9000 25.1000 48.2000 26.8000 ;
	    RECT 52.6000 26.8000 53.0000 27.2000 ;
	    RECT 54.2000 27.1000 54.5000 27.5000 ;
	    RECT 54.9000 27.4000 55.3000 27.5000 ;
	    RECT 56.6000 27.4000 57.0000 27.5000 ;
	    RECT 54.2000 26.8000 57.0000 27.1000 ;
	    RECT 52.6000 26.2000 52.9000 26.8000 ;
	    RECT 52.6000 25.8000 53.0000 26.2000 ;
	    RECT 44.7000 24.7000 45.1000 25.1000 ;
	    RECT 47.8000 24.7000 48.2000 25.1000 ;
	    RECT 54.2000 25.1000 54.5000 26.8000 ;
	    RECT 56.7000 26.1000 57.0000 26.8000 ;
	    RECT 56.7000 25.7000 57.1000 26.1000 ;
	    RECT 55.8000 25.1000 56.2000 25.2000 ;
	    RECT 56.6000 25.1000 57.0000 25.2000 ;
	    RECT 57.4000 25.1000 57.7000 27.5000 ;
	    RECT 54.2000 24.7000 54.6000 25.1000 ;
	    RECT 55.8000 24.8000 57.0000 25.1000 ;
	    RECT 57.3000 24.7000 57.7000 25.1000 ;
	    RECT 58.2000 26.8000 58.6000 27.2000 ;
	    RECT 42.2000 23.8000 42.6000 24.2000 ;
	    RECT 16.6000 22.8000 17.0000 23.2000 ;
	    RECT 16.6000 22.2000 16.9000 22.8000 ;
	    RECT 12.6000 21.8000 13.0000 22.2000 ;
	    RECT 15.0000 21.8000 15.4000 22.2000 ;
	    RECT 16.6000 21.8000 17.0000 22.2000 ;
	    RECT 9.4000 16.8000 9.8000 17.2000 ;
	    RECT 1.4000 15.9000 1.8000 16.3000 ;
	    RECT 4.5000 15.9000 4.9000 16.3000 ;
	    RECT 1.4000 14.2000 1.7000 15.9000 ;
	    RECT 3.9000 14.9000 4.3000 15.3000 ;
	    RECT 3.9000 14.2000 4.2000 14.9000 ;
	    RECT 1.4000 13.9000 4.2000 14.2000 ;
	    RECT 1.4000 13.5000 1.7000 13.9000 ;
	    RECT 2.1000 13.5000 2.5000 13.6000 ;
	    RECT 3.8000 13.5000 4.2000 13.6000 ;
	    RECT 4.6000 13.5000 4.9000 15.9000 ;
	    RECT 9.4000 16.2000 9.7000 16.8000 ;
	    RECT 9.4000 15.8000 9.8000 16.2000 ;
	    RECT 10.2000 16.1000 10.6000 16.2000 ;
	    RECT 11.0000 16.1000 11.4000 16.2000 ;
	    RECT 10.2000 15.8000 11.4000 16.1000 ;
	    RECT 7.0000 15.1000 7.4000 15.2000 ;
	    RECT 7.8000 15.1000 8.2000 15.2000 ;
	    RECT 7.0000 14.8000 8.2000 15.1000 ;
	    RECT 9.4000 14.8000 9.8000 15.2000 ;
	    RECT 9.4000 14.2000 9.7000 14.8000 ;
	    RECT 9.4000 14.1000 9.8000 14.2000 ;
	    RECT 10.2000 14.1000 10.6000 14.2000 ;
	    RECT 9.4000 13.8000 10.6000 14.1000 ;
	    RECT 11.8000 13.8000 12.2000 14.2000 ;
	    RECT 12.6000 14.1000 12.9000 21.8000 ;
	    RECT 13.4000 15.8000 13.8000 16.2000 ;
	    RECT 15.0000 16.1000 15.3000 21.8000 ;
	    RECT 29.4000 17.1000 29.8000 17.2000 ;
	    RECT 30.2000 17.1000 30.6000 17.2000 ;
	    RECT 29.4000 16.8000 30.6000 17.1000 ;
	    RECT 35.0000 16.8000 35.4000 17.2000 ;
	    RECT 41.4000 16.8000 41.8000 17.2000 ;
	    RECT 15.8000 16.1000 16.2000 16.2000 ;
	    RECT 15.0000 15.8000 16.2000 16.1000 ;
	    RECT 19.9000 15.9000 20.3000 16.3000 ;
	    RECT 23.0000 15.9000 23.4000 16.3000 ;
	    RECT 35.0000 16.2000 35.3000 16.8000 ;
	    RECT 41.4000 16.2000 41.7000 16.8000 ;
	    RECT 13.4000 15.2000 13.7000 15.8000 ;
	    RECT 13.4000 14.8000 13.8000 15.2000 ;
	    RECT 13.4000 14.1000 13.8000 14.2000 ;
	    RECT 12.6000 13.8000 13.8000 14.1000 ;
	    RECT 14.2000 13.8000 14.6000 14.2000 ;
	    RECT 15.8000 13.8000 16.2000 14.2000 ;
	    RECT 1.4000 13.1000 1.8000 13.5000 ;
	    RECT 2.1000 13.2000 4.9000 13.5000 ;
	    RECT 11.8000 13.2000 12.1000 13.8000 ;
	    RECT 4.5000 13.1000 4.9000 13.2000 ;
	    RECT 10.2000 12.8000 10.6000 13.2000 ;
	    RECT 11.8000 12.8000 12.2000 13.2000 ;
	    RECT 13.4000 13.1000 13.8000 13.2000 ;
	    RECT 14.2000 13.1000 14.5000 13.8000 ;
	    RECT 13.4000 12.8000 14.5000 13.1000 ;
	    RECT 3.0000 11.8000 3.4000 12.2000 ;
	    RECT 8.6000 11.8000 9.0000 12.2000 ;
	    RECT 3.0000 7.2000 3.3000 11.8000 ;
	    RECT 3.8000 7.5000 4.2000 7.9000 ;
	    RECT 6.9000 7.8000 7.3000 7.9000 ;
	    RECT 4.5000 7.5000 7.3000 7.8000 ;
	    RECT 3.0000 6.8000 3.4000 7.2000 ;
	    RECT 3.8000 7.1000 4.1000 7.5000 ;
	    RECT 4.5000 7.4000 4.9000 7.5000 ;
	    RECT 6.2000 7.4000 6.6000 7.5000 ;
	    RECT 3.8000 6.8000 6.6000 7.1000 ;
	    RECT 3.8000 5.1000 4.1000 6.8000 ;
	    RECT 6.3000 6.1000 6.6000 6.8000 ;
	    RECT 6.3000 5.7000 6.7000 6.1000 ;
	    RECT 7.0000 5.1000 7.3000 7.5000 ;
	    RECT 8.6000 7.2000 8.9000 11.8000 ;
	    RECT 8.6000 6.8000 9.0000 7.2000 ;
	    RECT 3.8000 4.7000 4.2000 5.1000 ;
	    RECT 6.9000 4.7000 7.3000 5.1000 ;
	    RECT 10.2000 6.2000 10.5000 12.8000 ;
	    RECT 11.0000 10.8000 11.4000 11.2000 ;
	    RECT 11.0000 9.2000 11.3000 10.8000 ;
	    RECT 11.0000 8.8000 11.4000 9.2000 ;
	    RECT 14.2000 8.2000 14.5000 12.8000 ;
	    RECT 15.0000 12.8000 15.4000 13.2000 ;
	    RECT 15.0000 12.2000 15.3000 12.8000 ;
	    RECT 15.0000 11.8000 15.4000 12.2000 ;
	    RECT 15.8000 11.2000 16.1000 13.8000 ;
	    RECT 19.9000 13.5000 20.2000 15.9000 ;
	    RECT 20.5000 14.9000 20.9000 15.3000 ;
	    RECT 20.6000 14.2000 20.9000 14.9000 ;
	    RECT 23.1000 14.2000 23.4000 15.9000 ;
	    RECT 27.0000 16.1000 27.4000 16.2000 ;
	    RECT 27.8000 16.1000 28.2000 16.2000 ;
	    RECT 27.0000 15.8000 28.2000 16.1000 ;
	    RECT 28.6000 15.8000 29.0000 16.2000 ;
	    RECT 31.0000 15.8000 31.4000 16.2000 ;
	    RECT 35.0000 15.8000 35.4000 16.2000 ;
	    RECT 38.2000 16.1000 38.6000 16.2000 ;
	    RECT 39.0000 16.1000 39.4000 16.2000 ;
	    RECT 38.2000 15.8000 39.4000 16.1000 ;
	    RECT 41.4000 15.8000 41.8000 16.2000 ;
	    RECT 20.6000 13.9000 23.4000 14.2000 ;
	    RECT 20.6000 13.5000 21.0000 13.6000 ;
	    RECT 22.3000 13.5000 22.7000 13.6000 ;
	    RECT 23.1000 13.5000 23.4000 13.9000 ;
	    RECT 19.9000 13.2000 22.7000 13.5000 ;
	    RECT 19.9000 13.1000 20.3000 13.2000 ;
	    RECT 23.0000 13.1000 23.4000 13.5000 ;
	    RECT 23.8000 13.8000 24.2000 14.2000 ;
	    RECT 27.0000 13.8000 27.4000 14.2000 ;
	    RECT 15.8000 10.8000 16.2000 11.2000 ;
	    RECT 23.8000 9.2000 24.1000 13.8000 ;
	    RECT 27.0000 12.2000 27.3000 13.8000 ;
	    RECT 27.0000 11.8000 27.4000 12.2000 ;
	    RECT 28.6000 9.2000 28.9000 15.8000 ;
	    RECT 29.4000 13.8000 29.8000 14.2000 ;
	    RECT 29.4000 13.2000 29.7000 13.8000 ;
	    RECT 29.4000 12.8000 29.8000 13.2000 ;
	    RECT 31.0000 9.2000 31.3000 15.8000 ;
	    RECT 39.8000 14.1000 40.2000 14.2000 ;
	    RECT 40.6000 14.1000 41.0000 14.2000 ;
	    RECT 39.8000 13.8000 41.0000 14.1000 ;
	    RECT 42.2000 13.2000 42.5000 23.8000 ;
	    RECT 50.2000 21.8000 50.6000 22.2000 ;
	    RECT 48.6000 17.1000 49.0000 17.2000 ;
	    RECT 49.4000 17.1000 49.8000 17.2000 ;
	    RECT 48.6000 16.8000 49.8000 17.1000 ;
	    RECT 50.2000 16.2000 50.5000 21.8000 ;
	    RECT 58.2000 19.2000 58.5000 26.8000 ;
	    RECT 59.0000 25.8000 59.4000 26.2000 ;
	    RECT 61.4000 25.8000 61.8000 26.2000 ;
	    RECT 59.0000 25.2000 59.3000 25.8000 ;
	    RECT 59.0000 24.8000 59.4000 25.2000 ;
	    RECT 61.4000 19.2000 61.7000 25.8000 ;
	    RECT 55.0000 19.1000 55.4000 19.2000 ;
	    RECT 55.8000 19.1000 56.2000 19.2000 ;
	    RECT 55.0000 18.8000 56.2000 19.1000 ;
	    RECT 58.2000 18.8000 58.6000 19.2000 ;
	    RECT 61.4000 18.8000 61.8000 19.2000 ;
	    RECT 43.8000 15.8000 44.2000 16.2000 ;
	    RECT 46.2000 16.1000 46.6000 16.2000 ;
	    RECT 47.0000 16.1000 47.4000 16.2000 ;
	    RECT 46.2000 15.8000 47.4000 16.1000 ;
	    RECT 50.2000 15.8000 50.6000 16.2000 ;
	    RECT 56.6000 15.8000 57.0000 16.2000 ;
	    RECT 59.9000 15.9000 60.3000 16.3000 ;
	    RECT 63.0000 15.9000 63.4000 16.3000 ;
	    RECT 43.8000 15.2000 44.1000 15.8000 ;
	    RECT 56.6000 15.2000 56.9000 15.8000 ;
	    RECT 43.8000 14.8000 44.2000 15.2000 ;
	    RECT 51.0000 15.1000 51.4000 15.2000 ;
	    RECT 51.8000 15.1000 52.2000 15.2000 ;
	    RECT 51.0000 14.8000 52.2000 15.1000 ;
	    RECT 56.6000 14.8000 57.0000 15.2000 ;
	    RECT 58.2000 14.8000 58.6000 15.2000 ;
	    RECT 43.8000 13.8000 44.2000 14.2000 ;
	    RECT 43.8000 13.2000 44.1000 13.8000 ;
	    RECT 32.6000 12.8000 33.0000 13.2000 ;
	    RECT 42.2000 12.8000 42.6000 13.2000 ;
	    RECT 43.8000 12.8000 44.2000 13.2000 ;
	    RECT 45.4000 13.1000 45.8000 13.2000 ;
	    RECT 44.6000 12.8000 45.8000 13.1000 ;
	    RECT 32.6000 9.2000 32.9000 12.8000 ;
	    RECT 40.6000 11.8000 41.0000 12.2000 ;
	    RECT 43.0000 12.1000 43.4000 12.2000 ;
	    RECT 43.0000 11.8000 44.1000 12.1000 ;
	    RECT 19.8000 9.1000 20.2000 9.2000 ;
	    RECT 20.6000 9.1000 21.0000 9.2000 ;
	    RECT 19.8000 8.8000 21.0000 9.1000 ;
	    RECT 23.8000 8.8000 24.2000 9.2000 ;
	    RECT 28.6000 8.8000 29.0000 9.2000 ;
	    RECT 31.0000 8.8000 31.4000 9.2000 ;
	    RECT 32.6000 8.8000 33.0000 9.2000 ;
	    RECT 31.0000 8.2000 31.3000 8.8000 ;
	    RECT 14.2000 7.8000 14.6000 8.2000 ;
	    RECT 18.2000 7.5000 18.6000 7.9000 ;
	    RECT 21.3000 7.8000 21.7000 7.9000 ;
	    RECT 18.9000 7.5000 21.7000 7.8000 ;
	    RECT 18.2000 7.1000 18.5000 7.5000 ;
	    RECT 18.9000 7.4000 19.3000 7.5000 ;
	    RECT 20.6000 7.4000 21.0000 7.5000 ;
	    RECT 18.2000 6.8000 21.0000 7.1000 ;
	    RECT 10.2000 5.8000 10.6000 6.2000 ;
	    RECT 10.2000 5.2000 10.5000 5.8000 ;
	    RECT 10.2000 4.8000 10.6000 5.2000 ;
	    RECT 18.2000 5.1000 18.5000 6.8000 ;
	    RECT 20.7000 6.1000 21.0000 6.8000 ;
	    RECT 20.7000 5.7000 21.1000 6.1000 ;
	    RECT 21.4000 5.1000 21.7000 7.5000 ;
	    RECT 26.2000 7.8000 26.6000 8.2000 ;
	    RECT 31.0000 7.8000 31.4000 8.2000 ;
	    RECT 31.8000 7.8000 32.2000 8.2000 ;
	    RECT 26.2000 7.2000 26.5000 7.8000 ;
	    RECT 31.8000 7.2000 32.1000 7.8000 ;
	    RECT 24.6000 7.1000 25.0000 7.2000 ;
	    RECT 25.4000 7.1000 25.8000 7.2000 ;
	    RECT 24.6000 6.8000 25.8000 7.1000 ;
	    RECT 26.2000 6.8000 26.6000 7.2000 ;
	    RECT 29.4000 7.1000 29.8000 7.2000 ;
	    RECT 30.2000 7.1000 30.6000 7.2000 ;
	    RECT 29.4000 6.8000 30.6000 7.1000 ;
	    RECT 31.8000 6.8000 32.2000 7.2000 ;
	    RECT 40.6000 6.2000 40.9000 11.8000 ;
	    RECT 43.8000 8.2000 44.1000 11.8000 ;
	    RECT 43.8000 7.8000 44.2000 8.2000 ;
	    RECT 18.2000 4.7000 18.6000 5.1000 ;
	    RECT 21.3000 4.7000 21.7000 5.1000 ;
	    RECT 24.6000 5.8000 25.0000 6.2000 ;
	    RECT 26.2000 6.1000 26.6000 6.2000 ;
	    RECT 27.0000 6.1000 27.4000 6.2000 ;
	    RECT 26.2000 5.8000 27.4000 6.1000 ;
	    RECT 33.4000 5.8000 33.8000 6.2000 ;
	    RECT 36.6000 5.8000 37.0000 6.2000 ;
	    RECT 40.6000 5.8000 41.0000 6.2000 ;
	    RECT 24.6000 5.2000 24.9000 5.8000 ;
	    RECT 33.4000 5.2000 33.7000 5.8000 ;
	    RECT 36.6000 5.2000 36.9000 5.8000 ;
	    RECT 44.6000 5.2000 44.9000 12.8000 ;
	    RECT 51.0000 9.1000 51.3000 14.8000 ;
	    RECT 58.2000 14.2000 58.5000 14.8000 ;
	    RECT 51.8000 13.8000 52.2000 14.2000 ;
	    RECT 58.2000 13.8000 58.6000 14.2000 ;
	    RECT 51.8000 13.2000 52.1000 13.8000 ;
	    RECT 59.9000 13.5000 60.2000 15.9000 ;
	    RECT 60.5000 14.9000 60.9000 15.3000 ;
	    RECT 60.6000 14.2000 60.9000 14.9000 ;
	    RECT 63.1000 14.2000 63.4000 15.9000 ;
	    RECT 60.6000 13.9000 63.4000 14.2000 ;
	    RECT 60.6000 13.5000 61.0000 13.6000 ;
	    RECT 62.3000 13.5000 62.7000 13.6000 ;
	    RECT 63.1000 13.5000 63.4000 13.9000 ;
	    RECT 59.9000 13.2000 62.7000 13.5000 ;
	    RECT 51.8000 12.8000 52.2000 13.2000 ;
	    RECT 52.6000 12.8000 53.0000 13.2000 ;
	    RECT 59.9000 13.1000 60.3000 13.2000 ;
	    RECT 63.0000 13.1000 63.4000 13.5000 ;
	    RECT 63.8000 13.8000 64.2000 14.2000 ;
	    RECT 51.8000 9.1000 52.2000 9.2000 ;
	    RECT 51.0000 8.8000 52.2000 9.1000 ;
	    RECT 49.4000 7.8000 49.8000 8.2000 ;
	    RECT 52.6000 8.1000 52.9000 12.8000 ;
	    RECT 63.8000 9.2000 64.1000 13.8000 ;
	    RECT 59.8000 9.1000 60.2000 9.2000 ;
	    RECT 60.6000 9.1000 61.0000 9.2000 ;
	    RECT 59.8000 8.8000 61.0000 9.1000 ;
	    RECT 63.8000 8.8000 64.2000 9.2000 ;
	    RECT 51.8000 7.8000 52.9000 8.1000 ;
	    RECT 49.4000 7.2000 49.7000 7.8000 ;
	    RECT 51.8000 7.2000 52.1000 7.8000 ;
	    RECT 58.2000 7.5000 58.6000 7.9000 ;
	    RECT 61.3000 7.8000 61.7000 7.9000 ;
	    RECT 58.9000 7.5000 61.7000 7.8000 ;
	    RECT 49.4000 6.8000 49.8000 7.2000 ;
	    RECT 51.8000 6.8000 52.2000 7.2000 ;
	    RECT 52.6000 7.1000 53.0000 7.2000 ;
	    RECT 53.4000 7.1000 53.8000 7.2000 ;
	    RECT 52.6000 6.8000 53.8000 7.1000 ;
	    RECT 58.2000 7.1000 58.5000 7.5000 ;
	    RECT 58.9000 7.4000 59.3000 7.5000 ;
	    RECT 60.6000 7.4000 61.0000 7.5000 ;
	    RECT 58.2000 6.8000 61.0000 7.1000 ;
	    RECT 53.4000 6.2000 53.7000 6.8000 ;
	    RECT 53.4000 5.8000 53.8000 6.2000 ;
	    RECT 54.2000 6.1000 54.6000 6.2000 ;
	    RECT 55.0000 6.1000 55.4000 6.2000 ;
	    RECT 54.2000 5.8000 55.4000 6.1000 ;
	    RECT 24.6000 4.8000 25.0000 5.2000 ;
	    RECT 30.2000 5.1000 30.6000 5.2000 ;
	    RECT 31.0000 5.1000 31.4000 5.2000 ;
	    RECT 30.2000 4.8000 31.4000 5.1000 ;
	    RECT 33.4000 4.8000 33.8000 5.2000 ;
	    RECT 36.6000 4.8000 37.0000 5.2000 ;
	    RECT 40.6000 5.1000 41.0000 5.2000 ;
	    RECT 41.4000 5.1000 41.8000 5.2000 ;
	    RECT 40.6000 4.8000 41.8000 5.1000 ;
	    RECT 44.6000 4.8000 45.0000 5.2000 ;
	    RECT 45.4000 5.1000 45.8000 5.2000 ;
	    RECT 46.2000 5.1000 46.6000 5.2000 ;
	    RECT 45.4000 4.8000 46.6000 5.1000 ;
	    RECT 51.8000 5.1000 52.2000 5.2000 ;
	    RECT 52.6000 5.1000 53.0000 5.2000 ;
	    RECT 51.8000 4.8000 53.0000 5.1000 ;
	    RECT 53.4000 4.8000 53.8000 5.2000 ;
	    RECT 58.2000 5.1000 58.5000 6.8000 ;
	    RECT 60.7000 6.1000 61.0000 6.8000 ;
	    RECT 60.7000 5.7000 61.1000 6.1000 ;
	    RECT 61.4000 5.1000 61.7000 7.5000 ;
	    RECT 53.4000 4.2000 53.7000 4.8000 ;
	    RECT 58.2000 4.7000 58.6000 5.1000 ;
	    RECT 61.3000 4.7000 61.7000 5.1000 ;
	    RECT 53.4000 3.8000 53.8000 4.2000 ;
         LAYER metal3 ;
	    RECT 32.6000 28.8000 33.0000 29.2000 ;
	    RECT 1.4000 27.8000 1.8000 28.2000 ;
	    RECT 31.0000 28.1000 31.4000 28.2000 ;
	    RECT 32.6000 28.1000 32.9000 28.8000 ;
	    RECT 30.2000 27.8000 32.9000 28.1000 ;
	    RECT 1.4000 27.1000 1.7000 27.8000 ;
	    RECT 11.0000 27.1000 11.4000 27.2000 ;
	    RECT 12.6000 27.1000 13.0000 27.2000 ;
	    RECT 1.4000 26.8000 13.0000 27.1000 ;
	    RECT 18.2000 27.1000 18.6000 27.2000 ;
	    RECT 25.4000 27.1000 25.8000 27.2000 ;
	    RECT 28.6000 27.1000 29.0000 27.2000 ;
	    RECT 18.2000 26.8000 29.0000 27.1000 ;
	    RECT 5.4000 26.1000 5.8000 26.2000 ;
	    RECT 19.0000 26.1000 19.4000 26.2000 ;
	    RECT 5.4000 25.8000 19.4000 26.1000 ;
	    RECT 29.4000 26.1000 29.8000 26.2000 ;
	    RECT 30.2000 26.1000 30.6000 26.2000 ;
	    RECT 29.4000 25.8000 30.6000 26.1000 ;
	    RECT 35.8000 26.1000 36.2000 26.2000 ;
	    RECT 39.8000 26.1000 40.2000 26.2000 ;
	    RECT 35.8000 25.8000 40.2000 26.1000 ;
	    RECT 47.0000 26.1000 47.4000 26.2000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 47.0000 25.8000 53.0000 26.1000 ;
	    RECT 9.4000 25.1000 9.8000 25.2000 ;
	    RECT 14.2000 25.1000 14.6000 25.2000 ;
	    RECT 9.4000 24.8000 14.6000 25.1000 ;
	    RECT 23.0000 25.1000 23.4000 25.2000 ;
	    RECT 26.2000 25.1000 26.6000 25.2000 ;
	    RECT 23.0000 24.8000 26.6000 25.1000 ;
	    RECT 55.8000 25.1000 56.2000 25.2000 ;
	    RECT 59.0000 25.1000 59.4000 25.2000 ;
	    RECT 55.8000 24.8000 59.4000 25.1000 ;
	    RECT 16.6000 22.8000 17.0000 23.2000 ;
	    RECT 15.0000 22.1000 15.4000 22.2000 ;
	    RECT 16.6000 22.1000 16.9000 22.8000 ;
	    RECT 15.0000 21.8000 16.9000 22.1000 ;
	    RECT 55.8000 19.1000 56.2000 19.2000 ;
	    RECT 58.2000 19.1000 58.6000 19.2000 ;
	    RECT 55.8000 18.8000 58.6000 19.1000 ;
	    RECT 30.2000 17.1000 30.6000 17.2000 ;
	    RECT 35.0000 17.1000 35.4000 17.2000 ;
	    RECT 48.6000 17.1000 49.0000 17.2000 ;
	    RECT 30.2000 16.8000 35.4000 17.1000 ;
	    RECT 41.4000 16.8000 49.0000 17.1000 ;
	    RECT 41.4000 16.2000 41.7000 16.8000 ;
	    RECT 9.4000 16.1000 9.8000 16.2000 ;
	    RECT 10.2000 16.1000 10.6000 16.2000 ;
	    RECT 13.4000 16.1000 13.8000 16.2000 ;
	    RECT 9.4000 15.8000 13.8000 16.1000 ;
	    RECT 27.8000 16.1000 28.2000 16.2000 ;
	    RECT 38.2000 16.1000 38.6000 16.2000 ;
	    RECT 27.8000 15.8000 38.6000 16.1000 ;
	    RECT 41.4000 15.8000 41.8000 16.2000 ;
	    RECT 43.8000 16.1000 44.2000 16.2000 ;
	    RECT 47.0000 16.1000 47.4000 16.2000 ;
	    RECT 50.2000 16.1000 50.6000 16.2000 ;
	    RECT 43.8000 15.8000 50.6000 16.1000 ;
	    RECT 7.8000 15.1000 8.2000 15.2000 ;
	    RECT 9.4000 15.1000 9.8000 15.2000 ;
	    RECT 7.8000 14.8000 9.8000 15.1000 ;
	    RECT 51.8000 15.1000 52.2000 15.2000 ;
	    RECT 56.6000 15.1000 57.0000 15.2000 ;
	    RECT 51.8000 14.8000 57.0000 15.1000 ;
	    RECT 10.2000 14.1000 10.6000 14.2000 ;
	    RECT 11.8000 14.1000 12.2000 14.2000 ;
	    RECT 10.2000 13.8000 12.2000 14.1000 ;
	    RECT 14.2000 14.1000 14.6000 14.2000 ;
	    RECT 40.6000 14.1000 41.0000 14.2000 ;
	    RECT 58.2000 14.1000 58.6000 14.2000 ;
	    RECT 14.2000 13.8000 29.7000 14.1000 ;
	    RECT 40.6000 13.8000 58.6000 14.1000 ;
	    RECT 29.4000 13.2000 29.7000 13.8000 ;
	    RECT 29.4000 12.8000 29.8000 13.2000 ;
	    RECT 42.2000 13.1000 42.6000 13.2000 ;
	    RECT 43.8000 13.1000 44.2000 13.2000 ;
	    RECT 42.2000 12.8000 44.2000 13.1000 ;
	    RECT 45.4000 13.1000 45.8000 13.2000 ;
	    RECT 51.8000 13.1000 52.2000 13.2000 ;
	    RECT 45.4000 12.8000 52.2000 13.1000 ;
	    RECT 8.6000 12.1000 9.0000 12.2000 ;
	    RECT 15.0000 12.1000 15.4000 12.2000 ;
	    RECT 27.0000 12.1000 27.4000 12.2000 ;
	    RECT 8.6000 11.8000 27.4000 12.1000 ;
	    RECT 11.0000 11.1000 11.4000 11.2000 ;
	    RECT 15.8000 11.1000 16.2000 11.2000 ;
	    RECT 11.0000 10.8000 16.2000 11.1000 ;
	    RECT 20.6000 9.1000 21.0000 9.2000 ;
	    RECT 23.8000 9.1000 24.2000 9.2000 ;
	    RECT 20.6000 8.8000 24.2000 9.1000 ;
	    RECT 60.6000 9.1000 61.0000 9.2000 ;
	    RECT 63.8000 9.1000 64.2000 9.2000 ;
	    RECT 60.6000 8.8000 64.2000 9.1000 ;
	    RECT 26.2000 8.1000 26.6000 8.2000 ;
	    RECT 31.0000 8.1000 31.4000 8.2000 ;
	    RECT 26.2000 7.8000 31.4000 8.1000 ;
	    RECT 24.6000 7.1000 25.0000 7.2000 ;
	    RECT 30.2000 7.1000 30.6000 7.2000 ;
	    RECT 31.8000 7.1000 32.2000 7.2000 ;
	    RECT 24.6000 6.8000 32.2000 7.1000 ;
	    RECT 49.4000 7.1000 49.8000 7.2000 ;
	    RECT 52.6000 7.1000 53.0000 7.2000 ;
	    RECT 49.4000 6.8000 53.0000 7.1000 ;
	    RECT 10.2000 6.1000 10.6000 6.2000 ;
	    RECT 26.2000 6.1000 26.6000 6.2000 ;
	    RECT 10.2000 5.8000 26.6000 6.1000 ;
	    RECT 36.6000 6.1000 37.0000 6.2000 ;
	    RECT 40.6000 6.1000 41.0000 6.2000 ;
	    RECT 36.6000 5.8000 41.0000 6.1000 ;
	    RECT 53.4000 6.1000 53.8000 6.2000 ;
	    RECT 54.2000 6.1000 54.6000 6.2000 ;
	    RECT 53.4000 5.8000 54.6000 6.1000 ;
	    RECT 24.6000 5.1000 25.0000 5.2000 ;
	    RECT 30.2000 5.1000 30.6000 5.2000 ;
	    RECT 33.4000 5.1000 33.8000 5.2000 ;
	    RECT 24.6000 4.8000 33.8000 5.1000 ;
	    RECT 41.4000 5.1000 41.8000 5.2000 ;
	    RECT 45.4000 5.1000 45.8000 5.2000 ;
	    RECT 41.4000 4.8000 45.8000 5.1000 ;
	    RECT 52.6000 5.1000 53.0000 5.2000 ;
	    RECT 53.4000 5.1000 53.8000 5.2000 ;
	    RECT 52.6000 4.8000 53.8000 5.1000 ;
   END
END adder
